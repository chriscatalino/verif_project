
module CannyEdge_DW01_addsub_1 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign B_AS[31] = B[31];
  assign B_AS[30] = B[30];
  assign B_AS[29] = B[29];
  assign B_AS[28] = B[28];
  assign B_AS[27] = B[27];
  assign B_AS[26] = B[26];
  assign B_AS[25] = B[25];
  assign B_AS[24] = B[24];
  assign B_AS[23] = B[23];
  assign B_AS[22] = B[22];
  assign B_AS[21] = B[21];
  assign B_AS[20] = B[20];
  assign B_AS[19] = B[19];
  assign B_AS[18] = B[18];
  assign B_AS[17] = B[17];
  assign B_AS[16] = B[16];
  assign B_AS[15] = B[15];
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_addsub_3 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n24,
         n25, n26, n27, n28, n29, n30;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];

  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  OAI21X1 U10 ( .A(n10), .B(n28), .C(n11), .Y(carry[7]) );
  OAI21X1 U11 ( .A(A[6]), .B(n22), .C(B[6]), .Y(n11) );
  AOI21X1 U12 ( .A(n12), .B(A[5]), .C(n23), .Y(n10) );
  OAI21X1 U13 ( .A(A[5]), .B(n12), .C(B[5]), .Y(n13) );
  OAI21X1 U14 ( .A(n14), .B(n29), .C(n15), .Y(n12) );
  OAI21X1 U15 ( .A(A[4]), .B(n24), .C(B[4]), .Y(n15) );
  AOI21X1 U16 ( .A(n16), .B(A[3]), .C(n25), .Y(n14) );
  OAI21X1 U17 ( .A(A[3]), .B(n16), .C(B[3]), .Y(n17) );
  OAI21X1 U18 ( .A(n18), .B(n30), .C(n19), .Y(n16) );
  OAI21X1 U19 ( .A(A[2]), .B(n26), .C(B[2]), .Y(n19) );
  AOI22X1 U20 ( .A(A[1]), .B(B[1]), .C(B[0]), .D(n27), .Y(n18) );
  OAI21X1 U21 ( .A(A[1]), .B(B[1]), .C(A[0]), .Y(n20) );
  INVX2 U1 ( .A(n10), .Y(n22) );
  INVX2 U2 ( .A(n13), .Y(n23) );
  INVX2 U3 ( .A(n14), .Y(n24) );
  INVX2 U4 ( .A(n17), .Y(n25) );
  INVX2 U5 ( .A(n18), .Y(n26) );
  INVX2 U6 ( .A(n20), .Y(n27) );
  INVX2 U7 ( .A(A[6]), .Y(n28) );
  INVX2 U8 ( .A(A[4]), .Y(n29) );
  INVX2 U9 ( .A(A[2]), .Y(n30) );
endmodule


module CannyEdge_DW01_addsub_4 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_0 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[0] = B[0];

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_1 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_2 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[0] = A[0];
  assign SUM[14] = carry[14];

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_4 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_7 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_8 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_9 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[14] = carry[14];

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_10 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_11 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_12 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n16), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n9), .B(B[28]), .Y(n1) );
  AND2X2 U2 ( .A(n10), .B(B[26]), .Y(n2) );
  AND2X2 U3 ( .A(n11), .B(B[24]), .Y(n3) );
  AND2X2 U4 ( .A(n12), .B(B[22]), .Y(n4) );
  AND2X2 U5 ( .A(n13), .B(B[20]), .Y(n5) );
  AND2X2 U6 ( .A(n14), .B(B[18]), .Y(n6) );
  AND2X2 U7 ( .A(n15), .B(B[16]), .Y(n7) );
  AND2X2 U8 ( .A(n1), .B(B[29]), .Y(n8) );
  AND2X2 U9 ( .A(n2), .B(B[27]), .Y(n9) );
  AND2X2 U10 ( .A(n3), .B(B[25]), .Y(n10) );
  AND2X2 U11 ( .A(n4), .B(B[23]), .Y(n11) );
  AND2X2 U12 ( .A(n5), .B(B[21]), .Y(n12) );
  AND2X2 U13 ( .A(n6), .B(B[19]), .Y(n13) );
  AND2X2 U14 ( .A(n7), .B(B[17]), .Y(n14) );
  AND2X2 U15 ( .A(carry[15]), .B(B[15]), .Y(n15) );
  AND2X2 U16 ( .A(B[0]), .B(A[0]), .Y(n16) );
  AND2X2 U17 ( .A(n8), .B(B[30]), .Y(n17) );
  XOR2X1 U18 ( .A(B[31]), .B(n17), .Y(SUM[31]) );
  XOR2X1 U19 ( .A(n8), .B(B[30]), .Y(SUM[30]) );
  XOR2X1 U20 ( .A(n1), .B(B[29]), .Y(SUM[29]) );
  XOR2X1 U21 ( .A(n9), .B(B[28]), .Y(SUM[28]) );
  XOR2X1 U22 ( .A(n2), .B(B[27]), .Y(SUM[27]) );
  XOR2X1 U23 ( .A(n10), .B(B[26]), .Y(SUM[26]) );
  XOR2X1 U24 ( .A(n3), .B(B[25]), .Y(SUM[25]) );
  XOR2X1 U25 ( .A(n11), .B(B[24]), .Y(SUM[24]) );
  XOR2X1 U26 ( .A(n4), .B(B[23]), .Y(SUM[23]) );
  XOR2X1 U27 ( .A(n12), .B(B[22]), .Y(SUM[22]) );
  XOR2X1 U28 ( .A(n5), .B(B[21]), .Y(SUM[21]) );
  XOR2X1 U29 ( .A(n13), .B(B[20]), .Y(SUM[20]) );
  XOR2X1 U30 ( .A(n6), .B(B[19]), .Y(SUM[19]) );
  XOR2X1 U31 ( .A(n14), .B(B[18]), .Y(SUM[18]) );
  XOR2X1 U32 ( .A(n7), .B(B[17]), .Y(SUM[17]) );
  XOR2X1 U33 ( .A(n15), .B(B[16]), .Y(SUM[16]) );
  XOR2X1 U34 ( .A(carry[15]), .B(B[15]), .Y(SUM[15]) );
  XOR2X1 U35 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_13 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1;
  wire   [9:1] carry;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U2 ( .A(carry[8]), .B(B[8]), .Y(SUM[9]) );
  XOR2X1 U3 ( .A(carry[8]), .B(B[8]), .Y(SUM[8]) );
  XOR2X1 U4 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_14 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n8), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n10), .B(A[28]), .Y(n1) );
  AND2X2 U2 ( .A(n11), .B(A[26]), .Y(n2) );
  AND2X2 U3 ( .A(n12), .B(A[24]), .Y(n3) );
  AND2X2 U4 ( .A(n13), .B(A[22]), .Y(n4) );
  AND2X2 U5 ( .A(n14), .B(A[20]), .Y(n5) );
  AND2X2 U6 ( .A(n15), .B(A[18]), .Y(n6) );
  AND2X2 U7 ( .A(n16), .B(A[16]), .Y(n7) );
  AND2X2 U8 ( .A(B[0]), .B(A[0]), .Y(n8) );
  AND2X2 U9 ( .A(n1), .B(A[29]), .Y(n9) );
  AND2X2 U10 ( .A(n2), .B(A[27]), .Y(n10) );
  AND2X2 U11 ( .A(n3), .B(A[25]), .Y(n11) );
  AND2X2 U12 ( .A(n4), .B(A[23]), .Y(n12) );
  AND2X2 U13 ( .A(n5), .B(A[21]), .Y(n13) );
  AND2X2 U14 ( .A(n6), .B(A[19]), .Y(n14) );
  AND2X2 U15 ( .A(n7), .B(A[17]), .Y(n15) );
  AND2X2 U16 ( .A(carry[15]), .B(A[15]), .Y(n16) );
  AND2X2 U17 ( .A(n9), .B(A[30]), .Y(n17) );
  XOR2X1 U18 ( .A(A[31]), .B(n17), .Y(SUM[31]) );
  XOR2X1 U19 ( .A(n9), .B(A[30]), .Y(SUM[30]) );
  XOR2X1 U20 ( .A(n1), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U21 ( .A(n10), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U22 ( .A(n2), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U23 ( .A(n11), .B(A[26]), .Y(SUM[26]) );
  XOR2X1 U24 ( .A(n3), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U25 ( .A(n12), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U26 ( .A(n4), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U27 ( .A(n13), .B(A[22]), .Y(SUM[22]) );
  XOR2X1 U28 ( .A(n5), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U29 ( .A(n14), .B(A[20]), .Y(SUM[20]) );
  XOR2X1 U30 ( .A(n6), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U31 ( .A(n15), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U32 ( .A(n7), .B(A[17]), .Y(SUM[17]) );
  XOR2X1 U33 ( .A(n16), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U34 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U35 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_15 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_16 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_17 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_18 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U3 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_addsub_5 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign SUM[0] = A[0];
  assign SUM[14] = carry[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];

  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B_AS[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_addsub_7 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  XOR2X1 U1 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[31]), .B(carry[0]), .Y(B_AS[31]) );
  XOR2X1 U9 ( .A(B[30]), .B(carry[0]), .Y(B_AS[30]) );
  XOR2X1 U10 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U11 ( .A(B[29]), .B(carry[0]), .Y(B_AS[29]) );
  XOR2X1 U12 ( .A(B[28]), .B(carry[0]), .Y(B_AS[28]) );
  XOR2X1 U13 ( .A(B[27]), .B(carry[0]), .Y(B_AS[27]) );
  XOR2X1 U14 ( .A(B[26]), .B(carry[0]), .Y(B_AS[26]) );
  XOR2X1 U15 ( .A(B[25]), .B(carry[0]), .Y(B_AS[25]) );
  XOR2X1 U16 ( .A(B[24]), .B(carry[0]), .Y(B_AS[24]) );
  XOR2X1 U17 ( .A(B[23]), .B(carry[0]), .Y(B_AS[23]) );
  XOR2X1 U18 ( .A(B[22]), .B(carry[0]), .Y(B_AS[22]) );
  XOR2X1 U19 ( .A(B[21]), .B(carry[0]), .Y(B_AS[21]) );
  XOR2X1 U20 ( .A(B[20]), .B(carry[0]), .Y(B_AS[20]) );
  XOR2X1 U21 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U22 ( .A(B[19]), .B(carry[0]), .Y(B_AS[19]) );
  XOR2X1 U23 ( .A(B[18]), .B(carry[0]), .Y(B_AS[18]) );
  XOR2X1 U24 ( .A(B[17]), .B(carry[0]), .Y(B_AS[17]) );
  XOR2X1 U25 ( .A(B[16]), .B(carry[0]), .Y(B_AS[16]) );
  XOR2X1 U26 ( .A(B[15]), .B(carry[0]), .Y(B_AS[15]) );
  XOR2X1 U27 ( .A(B[14]), .B(carry[0]), .Y(B_AS[14]) );
  XOR2X1 U28 ( .A(B[13]), .B(carry[0]), .Y(B_AS[13]) );
  XOR2X1 U29 ( .A(B[12]), .B(carry[0]), .Y(B_AS[12]) );
  XOR2X1 U30 ( .A(B[11]), .B(carry[0]), .Y(B_AS[11]) );
  XOR2X1 U31 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U32 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_add_19 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_20 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [31:1] carry;

  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n9), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n11), .B(B[28]), .Y(n1) );
  AND2X2 U2 ( .A(n12), .B(B[26]), .Y(n2) );
  AND2X2 U3 ( .A(n13), .B(B[24]), .Y(n3) );
  AND2X2 U4 ( .A(n14), .B(B[22]), .Y(n4) );
  AND2X2 U5 ( .A(n15), .B(B[20]), .Y(n5) );
  AND2X2 U6 ( .A(n16), .B(B[18]), .Y(n6) );
  AND2X2 U7 ( .A(n17), .B(B[16]), .Y(n7) );
  AND2X2 U8 ( .A(n22), .B(B[14]), .Y(n8) );
  AND2X2 U9 ( .A(B[0]), .B(A[0]), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(B[29]), .Y(n10) );
  AND2X2 U11 ( .A(n2), .B(B[27]), .Y(n11) );
  AND2X2 U12 ( .A(n3), .B(B[25]), .Y(n12) );
  AND2X2 U13 ( .A(n4), .B(B[23]), .Y(n13) );
  AND2X2 U14 ( .A(n5), .B(B[21]), .Y(n14) );
  AND2X2 U15 ( .A(n6), .B(B[19]), .Y(n15) );
  AND2X2 U16 ( .A(n7), .B(B[17]), .Y(n16) );
  AND2X2 U17 ( .A(n8), .B(B[15]), .Y(n17) );
  AND2X2 U18 ( .A(carry[9]), .B(B[9]), .Y(n18) );
  AND2X2 U19 ( .A(n18), .B(B[10]), .Y(n19) );
  AND2X2 U20 ( .A(n19), .B(B[11]), .Y(n20) );
  AND2X2 U21 ( .A(n20), .B(B[12]), .Y(n21) );
  AND2X2 U22 ( .A(n21), .B(B[13]), .Y(n22) );
  AND2X2 U23 ( .A(n10), .B(B[30]), .Y(n23) );
  XOR2X1 U24 ( .A(B[31]), .B(n23), .Y(SUM[31]) );
  XOR2X1 U25 ( .A(n10), .B(B[30]), .Y(SUM[30]) );
  XOR2X1 U26 ( .A(n1), .B(B[29]), .Y(SUM[29]) );
  XOR2X1 U27 ( .A(n11), .B(B[28]), .Y(SUM[28]) );
  XOR2X1 U28 ( .A(n2), .B(B[27]), .Y(SUM[27]) );
  XOR2X1 U29 ( .A(n12), .B(B[26]), .Y(SUM[26]) );
  XOR2X1 U30 ( .A(n3), .B(B[25]), .Y(SUM[25]) );
  XOR2X1 U31 ( .A(n13), .B(B[24]), .Y(SUM[24]) );
  XOR2X1 U32 ( .A(n4), .B(B[23]), .Y(SUM[23]) );
  XOR2X1 U33 ( .A(n14), .B(B[22]), .Y(SUM[22]) );
  XOR2X1 U34 ( .A(n5), .B(B[21]), .Y(SUM[21]) );
  XOR2X1 U35 ( .A(n15), .B(B[20]), .Y(SUM[20]) );
  XOR2X1 U36 ( .A(n6), .B(B[19]), .Y(SUM[19]) );
  XOR2X1 U37 ( .A(n16), .B(B[18]), .Y(SUM[18]) );
  XOR2X1 U38 ( .A(n7), .B(B[17]), .Y(SUM[17]) );
  XOR2X1 U39 ( .A(n17), .B(B[16]), .Y(SUM[16]) );
  XOR2X1 U40 ( .A(n8), .B(B[15]), .Y(SUM[15]) );
  XOR2X1 U41 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U42 ( .A(carry[9]), .B(B[9]), .Y(SUM[9]) );
  XOR2X1 U43 ( .A(n18), .B(B[10]), .Y(SUM[10]) );
  XOR2X1 U44 ( .A(n19), .B(B[11]), .Y(SUM[11]) );
  XOR2X1 U45 ( .A(n20), .B(B[12]), .Y(SUM[12]) );
  XOR2X1 U46 ( .A(n21), .B(B[13]), .Y(SUM[13]) );
  XOR2X1 U47 ( .A(n22), .B(B[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_add_21 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [31:1] carry;

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n9), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n10), .B(A[29]), .Y(n1) );
  AND2X2 U2 ( .A(n11), .B(A[27]), .Y(n2) );
  AND2X2 U3 ( .A(n12), .B(A[25]), .Y(n3) );
  AND2X2 U4 ( .A(n13), .B(A[23]), .Y(n4) );
  AND2X2 U5 ( .A(n14), .B(A[21]), .Y(n5) );
  AND2X2 U6 ( .A(n15), .B(A[19]), .Y(n6) );
  AND2X2 U7 ( .A(n16), .B(A[17]), .Y(n7) );
  AND2X2 U8 ( .A(n17), .B(A[15]), .Y(n8) );
  AND2X2 U9 ( .A(B[0]), .B(A[0]), .Y(n9) );
  AND2X2 U10 ( .A(n2), .B(A[28]), .Y(n10) );
  AND2X2 U11 ( .A(n3), .B(A[26]), .Y(n11) );
  AND2X2 U12 ( .A(n4), .B(A[24]), .Y(n12) );
  AND2X2 U13 ( .A(n5), .B(A[22]), .Y(n13) );
  AND2X2 U14 ( .A(n6), .B(A[20]), .Y(n14) );
  AND2X2 U15 ( .A(n7), .B(A[18]), .Y(n15) );
  AND2X2 U16 ( .A(n8), .B(A[16]), .Y(n16) );
  AND2X2 U17 ( .A(carry[14]), .B(A[14]), .Y(n17) );
  AND2X2 U18 ( .A(n1), .B(A[30]), .Y(n18) );
  XOR2X1 U19 ( .A(A[31]), .B(n18), .Y(SUM[31]) );
  XOR2X1 U20 ( .A(n1), .B(A[30]), .Y(SUM[30]) );
  XOR2X1 U21 ( .A(n10), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U22 ( .A(n2), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U23 ( .A(n11), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U24 ( .A(n3), .B(A[26]), .Y(SUM[26]) );
  XOR2X1 U25 ( .A(n12), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U26 ( .A(n4), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U27 ( .A(n13), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U28 ( .A(n5), .B(A[22]), .Y(SUM[22]) );
  XOR2X1 U29 ( .A(n14), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U30 ( .A(n6), .B(A[20]), .Y(SUM[20]) );
  XOR2X1 U31 ( .A(n15), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U32 ( .A(n7), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U33 ( .A(n16), .B(A[17]), .Y(SUM[17]) );
  XOR2X1 U34 ( .A(n8), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U35 ( .A(n17), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U36 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U37 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_addsub_9 ( A, B, CI, ADD_SUB, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [7:0] carry;
  wire   [6:0] B_AS;
  assign B_AS[6] = B[6];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[6]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[6]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_addsub_11 ( A, B, CI, ADD_SUB, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n12, n13, n14, n15;
  wire   [11:0] carry;
  wire   [10:0] B_AS;

  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YS(SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  OAI21X1 U5 ( .A(n12), .B(n15), .C(n5), .Y(carry[3]) );
  OAI21X1 U6 ( .A(A[2]), .B(n6), .C(n7), .Y(n5) );
  XOR2X1 U7 ( .A(B[2]), .B(ADD_SUB), .Y(n7) );
  OAI21X1 U8 ( .A(n8), .B(n14), .C(n9), .Y(n6) );
  OAI21X1 U9 ( .A(A[1]), .B(n13), .C(n10), .Y(n9) );
  XOR2X1 U10 ( .A(B[1]), .B(ADD_SUB), .Y(n10) );
  MUX2X1 U11 ( .B(ADD_SUB), .A(A[0]), .S(B[0]), .Y(n8) );
  XOR2X1 U12 ( .A(B[9]), .B(ADD_SUB), .Y(B_AS[9]) );
  XOR2X1 U13 ( .A(B[8]), .B(ADD_SUB), .Y(B_AS[8]) );
  XOR2X1 U14 ( .A(B[7]), .B(ADD_SUB), .Y(B_AS[7]) );
  XOR2X1 U15 ( .A(B[6]), .B(ADD_SUB), .Y(B_AS[6]) );
  XOR2X1 U16 ( .A(B[5]), .B(ADD_SUB), .Y(B_AS[5]) );
  XOR2X1 U17 ( .A(B[4]), .B(ADD_SUB), .Y(B_AS[4]) );
  XOR2X1 U18 ( .A(B[3]), .B(ADD_SUB), .Y(B_AS[3]) );
  XOR2X1 U19 ( .A(B[10]), .B(ADD_SUB), .Y(B_AS[10]) );
  INVX2 U1 ( .A(n6), .Y(n12) );
  INVX2 U2 ( .A(n8), .Y(n13) );
  INVX2 U3 ( .A(A[1]), .Y(n14) );
  INVX2 U4 ( .A(A[2]), .Y(n15) );
endmodule


module CannyEdge_DW01_addsub_12 ( A, B, CI, ADD_SUB, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [11:0] carry;
  wire   [10:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YS(SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  XOR2X1 U1 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U9 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U10 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U11 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;
  tri   [31:0] A;

  OAI21X1 U59 ( .A(B[31]), .B(n59), .C(n60), .Y(LT_LE) );
  OAI21X1 U60 ( .A(n135), .B(n61), .C(A[31]), .Y(n60) );
  NAND2X1 U61 ( .A(A[30]), .B(n59), .Y(n61) );
  OAI21X1 U62 ( .A(B[31]), .B(n177), .C(n62), .Y(n59) );
  AOI21X1 U63 ( .A(A[29]), .B(n134), .C(n63), .Y(n62) );
  AOI21X1 U64 ( .A(B[29]), .B(n176), .C(n64), .Y(n63) );
  OAI21X1 U65 ( .A(A[28]), .B(n133), .C(n65), .Y(n64) );
  OAI21X1 U66 ( .A(B[28]), .B(n175), .C(n66), .Y(n65) );
  AOI21X1 U67 ( .A(A[27]), .B(n132), .C(n67), .Y(n66) );
  AOI21X1 U68 ( .A(B[27]), .B(n174), .C(n68), .Y(n67) );
  OAI21X1 U69 ( .A(A[26]), .B(n131), .C(n69), .Y(n68) );
  OAI21X1 U70 ( .A(B[26]), .B(n173), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(A[25]), .B(n130), .C(n71), .Y(n70) );
  AOI21X1 U72 ( .A(B[25]), .B(n172), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(A[24]), .B(n129), .C(n73), .Y(n72) );
  OAI21X1 U74 ( .A(B[24]), .B(n171), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(A[23]), .B(n128), .C(n75), .Y(n74) );
  AOI21X1 U76 ( .A(B[23]), .B(n170), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(A[22]), .B(n127), .C(n77), .Y(n76) );
  OAI21X1 U78 ( .A(B[22]), .B(n169), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(A[21]), .B(n126), .C(n79), .Y(n78) );
  AOI21X1 U80 ( .A(B[21]), .B(n168), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(A[20]), .B(n125), .C(n81), .Y(n80) );
  OAI21X1 U82 ( .A(B[20]), .B(n167), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(A[19]), .B(n124), .C(n83), .Y(n82) );
  AOI21X1 U84 ( .A(B[19]), .B(n166), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(A[18]), .B(n123), .C(n85), .Y(n84) );
  OAI21X1 U86 ( .A(B[18]), .B(n165), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(A[17]), .B(n122), .C(n87), .Y(n86) );
  AOI21X1 U88 ( .A(B[17]), .B(n164), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(A[16]), .B(n121), .C(n89), .Y(n88) );
  OAI21X1 U90 ( .A(B[16]), .B(n163), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(A[15]), .B(n120), .C(n91), .Y(n90) );
  AOI21X1 U92 ( .A(B[15]), .B(n162), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(A[14]), .B(n136), .C(n93), .Y(n92) );
  OAI21X1 U94 ( .A(B[14]), .B(n161), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(A[13]), .B(n137), .C(n95), .Y(n94) );
  AOI21X1 U96 ( .A(B[13]), .B(n160), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(A[12]), .B(n138), .C(n97), .Y(n96) );
  OAI21X1 U98 ( .A(B[12]), .B(n159), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(A[11]), .B(n139), .C(n99), .Y(n98) );
  AOI21X1 U100 ( .A(B[11]), .B(n158), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(A[10]), .B(n140), .C(n101), .Y(n100) );
  OAI21X1 U102 ( .A(B[9]), .B(n157), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(A[10]), .B(n140), .C(n103), .Y(n102) );
  AOI21X1 U104 ( .A(B[9]), .B(n157), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(A[8]), .B(n141), .C(n105), .Y(n104) );
  OAI21X1 U106 ( .A(B[8]), .B(n156), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(A[7]), .B(n142), .C(n107), .Y(n106) );
  AOI21X1 U108 ( .A(B[7]), .B(n155), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(A[6]), .B(n143), .C(n109), .Y(n108) );
  OAI21X1 U110 ( .A(B[6]), .B(n154), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(A[5]), .B(n144), .C(n111), .Y(n110) );
  AOI21X1 U112 ( .A(B[5]), .B(n153), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(A[4]), .B(n145), .C(n113), .Y(n112) );
  OAI21X1 U114 ( .A(B[4]), .B(n152), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(A[3]), .B(n146), .C(n115), .Y(n114) );
  AOI21X1 U116 ( .A(B[3]), .B(n151), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(A[2]), .B(n147), .C(n117), .Y(n116) );
  OAI21X1 U118 ( .A(B[2]), .B(n150), .C(n118), .Y(n117) );
  AOI22X1 U119 ( .A(n119), .B(A[0]), .C(A[1]), .D(n148), .Y(n118) );
  AOI21X1 U120 ( .A(B[1]), .B(n149), .C(B[0]), .Y(n119) );
  INVX2 U1 ( .A(B[15]), .Y(n120) );
  INVX2 U2 ( .A(B[16]), .Y(n121) );
  INVX2 U3 ( .A(B[17]), .Y(n122) );
  INVX2 U4 ( .A(B[18]), .Y(n123) );
  INVX2 U5 ( .A(B[19]), .Y(n124) );
  INVX2 U6 ( .A(B[20]), .Y(n125) );
  INVX2 U7 ( .A(B[21]), .Y(n126) );
  INVX2 U8 ( .A(B[22]), .Y(n127) );
  INVX2 U9 ( .A(B[23]), .Y(n128) );
  INVX2 U10 ( .A(B[24]), .Y(n129) );
  INVX2 U11 ( .A(B[25]), .Y(n130) );
  INVX2 U12 ( .A(B[26]), .Y(n131) );
  INVX2 U13 ( .A(B[27]), .Y(n132) );
  INVX2 U14 ( .A(B[28]), .Y(n133) );
  INVX2 U15 ( .A(B[29]), .Y(n134) );
  INVX2 U16 ( .A(B[31]), .Y(n135) );
  INVX2 U17 ( .A(B[14]), .Y(n136) );
  INVX2 U18 ( .A(B[13]), .Y(n137) );
  INVX2 U19 ( .A(B[12]), .Y(n138) );
  INVX2 U20 ( .A(B[11]), .Y(n139) );
  INVX2 U21 ( .A(B[10]), .Y(n140) );
  INVX2 U22 ( .A(B[8]), .Y(n141) );
  INVX2 U23 ( .A(B[7]), .Y(n142) );
  INVX2 U24 ( .A(B[6]), .Y(n143) );
  INVX2 U25 ( .A(B[5]), .Y(n144) );
  INVX2 U26 ( .A(B[4]), .Y(n145) );
  INVX2 U27 ( .A(B[3]), .Y(n146) );
  INVX2 U28 ( .A(B[2]), .Y(n147) );
  INVX2 U29 ( .A(B[1]), .Y(n148) );
  INVX2 U30 ( .A(A[1]), .Y(n149) );
  INVX2 U31 ( .A(A[2]), .Y(n150) );
  INVX2 U32 ( .A(A[3]), .Y(n151) );
  INVX2 U33 ( .A(A[4]), .Y(n152) );
  INVX2 U34 ( .A(A[5]), .Y(n153) );
  INVX2 U35 ( .A(A[6]), .Y(n154) );
  INVX2 U36 ( .A(A[7]), .Y(n155) );
  INVX2 U37 ( .A(A[8]), .Y(n156) );
  INVX2 U38 ( .A(A[9]), .Y(n157) );
  INVX2 U39 ( .A(A[11]), .Y(n158) );
  INVX2 U40 ( .A(A[12]), .Y(n159) );
  INVX2 U41 ( .A(A[13]), .Y(n160) );
  INVX2 U42 ( .A(A[14]), .Y(n161) );
  INVX2 U43 ( .A(A[15]), .Y(n162) );
  INVX2 U44 ( .A(A[16]), .Y(n163) );
  INVX2 U45 ( .A(A[17]), .Y(n164) );
  INVX2 U46 ( .A(A[18]), .Y(n165) );
  INVX2 U47 ( .A(A[19]), .Y(n166) );
  INVX2 U48 ( .A(A[20]), .Y(n167) );
  INVX2 U49 ( .A(A[21]), .Y(n168) );
  INVX2 U50 ( .A(A[22]), .Y(n169) );
  INVX2 U51 ( .A(A[23]), .Y(n170) );
  INVX2 U52 ( .A(A[24]), .Y(n171) );
  INVX2 U53 ( .A(A[25]), .Y(n172) );
  INVX2 U54 ( .A(A[26]), .Y(n173) );
  INVX2 U55 ( .A(A[27]), .Y(n174) );
  INVX2 U56 ( .A(A[28]), .Y(n175) );
  INVX2 U57 ( .A(A[29]), .Y(n176) );
  INVX2 U58 ( .A(A[30]), .Y(n177) );
endmodule


module CannyEdge_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182;
  tri   [31:0] B;

  OAI21X1 U61 ( .A(n124), .B(n61), .C(n62), .Y(LT_LE) );
  OAI21X1 U62 ( .A(n123), .B(n63), .C(n182), .Y(n62) );
  OAI21X1 U64 ( .A(B[30]), .B(n124), .C(n64), .Y(n61) );
  AOI21X1 U65 ( .A(A[29]), .B(n181), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n137), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n180), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n136), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n179), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n135), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n178), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n134), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n177), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n133), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n176), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n132), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n175), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n131), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n174), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n130), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n173), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n129), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n172), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n128), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n171), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n127), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n170), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n126), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n169), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n125), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n168), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n138), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n167), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n139), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n166), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n140), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n165), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n141), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n164), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n142), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n163), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n143), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n162), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n144), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n162), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n144), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n161), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n145), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n160), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n146), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n159), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n147), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n158), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n148), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n149), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n156), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n150), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n155), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n151), .C(n120), .Y(n119) );
  AOI21X1 U121 ( .A(A[1]), .B(n121), .C(n152), .Y(n120) );
  OAI21X1 U122 ( .A(n121), .B(A[1]), .C(n154), .Y(n122) );
  NAND2X1 U123 ( .A(B[0]), .B(n153), .Y(n121) );
  OR2X2 U63 ( .A(A[31]), .B(B[30]), .Y(n63) );
  INVX2 U1 ( .A(n61), .Y(n123) );
  INVX2 U2 ( .A(A[31]), .Y(n124) );
  INVX2 U3 ( .A(A[17]), .Y(n125) );
  INVX2 U4 ( .A(A[18]), .Y(n126) );
  INVX2 U5 ( .A(A[19]), .Y(n127) );
  INVX2 U6 ( .A(A[20]), .Y(n128) );
  INVX2 U7 ( .A(A[21]), .Y(n129) );
  INVX2 U8 ( .A(A[22]), .Y(n130) );
  INVX2 U9 ( .A(A[23]), .Y(n131) );
  INVX2 U10 ( .A(A[24]), .Y(n132) );
  INVX2 U11 ( .A(A[25]), .Y(n133) );
  INVX2 U12 ( .A(A[26]), .Y(n134) );
  INVX2 U13 ( .A(A[27]), .Y(n135) );
  INVX2 U14 ( .A(A[28]), .Y(n136) );
  INVX2 U15 ( .A(A[29]), .Y(n137) );
  INVX2 U16 ( .A(A[16]), .Y(n138) );
  INVX2 U17 ( .A(A[15]), .Y(n139) );
  INVX2 U18 ( .A(A[14]), .Y(n140) );
  INVX2 U19 ( .A(A[13]), .Y(n141) );
  INVX2 U20 ( .A(A[12]), .Y(n142) );
  INVX2 U21 ( .A(A[11]), .Y(n143) );
  INVX2 U22 ( .A(A[9]), .Y(n144) );
  INVX2 U23 ( .A(A[8]), .Y(n145) );
  INVX2 U24 ( .A(A[7]), .Y(n146) );
  INVX2 U25 ( .A(A[6]), .Y(n147) );
  INVX2 U26 ( .A(A[5]), .Y(n148) );
  INVX2 U27 ( .A(A[4]), .Y(n149) );
  INVX2 U28 ( .A(A[3]), .Y(n150) );
  INVX2 U29 ( .A(A[2]), .Y(n151) );
  INVX2 U30 ( .A(n122), .Y(n152) );
  INVX2 U31 ( .A(A[0]), .Y(n153) );
  INVX2 U32 ( .A(B[1]), .Y(n154) );
  INVX2 U33 ( .A(B[2]), .Y(n155) );
  INVX2 U34 ( .A(B[3]), .Y(n156) );
  INVX2 U35 ( .A(B[4]), .Y(n157) );
  INVX2 U36 ( .A(B[5]), .Y(n158) );
  INVX2 U37 ( .A(B[6]), .Y(n159) );
  INVX2 U38 ( .A(B[7]), .Y(n160) );
  INVX2 U39 ( .A(B[8]), .Y(n161) );
  INVX2 U40 ( .A(B[10]), .Y(n162) );
  INVX2 U41 ( .A(B[11]), .Y(n163) );
  INVX2 U42 ( .A(B[12]), .Y(n164) );
  INVX2 U43 ( .A(B[13]), .Y(n165) );
  INVX2 U44 ( .A(B[14]), .Y(n166) );
  INVX2 U45 ( .A(B[15]), .Y(n167) );
  INVX2 U46 ( .A(B[16]), .Y(n168) );
  INVX2 U47 ( .A(B[17]), .Y(n169) );
  INVX2 U48 ( .A(B[18]), .Y(n170) );
  INVX2 U49 ( .A(B[19]), .Y(n171) );
  INVX2 U50 ( .A(B[20]), .Y(n172) );
  INVX2 U51 ( .A(B[21]), .Y(n173) );
  INVX2 U52 ( .A(B[22]), .Y(n174) );
  INVX2 U53 ( .A(B[23]), .Y(n175) );
  INVX2 U54 ( .A(B[24]), .Y(n176) );
  INVX2 U55 ( .A(B[25]), .Y(n177) );
  INVX2 U56 ( .A(B[26]), .Y(n178) );
  INVX2 U57 ( .A(B[27]), .Y(n179) );
  INVX2 U58 ( .A(B[28]), .Y(n180) );
  INVX2 U59 ( .A(B[29]), .Y(n181) );
  INVX2 U60 ( .A(B[31]), .Y(n182) );
endmodule


module CannyEdge_DW01_cmp2_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182;
  tri   [31:0] B;

  OAI21X1 U61 ( .A(n139), .B(n61), .C(n62), .Y(LT_LE) );
  OAI21X1 U62 ( .A(n123), .B(n63), .C(n182), .Y(n62) );
  OAI21X1 U64 ( .A(B[30]), .B(n139), .C(n64), .Y(n61) );
  AOI21X1 U65 ( .A(A[29]), .B(n181), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n138), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n180), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n137), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n179), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n136), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n178), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n135), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n177), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n134), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n176), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n133), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n175), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n132), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n174), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n131), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n173), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n130), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n172), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n129), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n171), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n128), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n170), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n127), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n169), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n126), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n168), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n125), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n167), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n124), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n166), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n140), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n165), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n141), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n164), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n142), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n163), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n143), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n162), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n144), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n162), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n144), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n161), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n145), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n160), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n146), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n159), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n147), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n158), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n148), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n149), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n156), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n150), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n155), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n151), .C(n120), .Y(n119) );
  AOI21X1 U121 ( .A(A[1]), .B(n121), .C(n152), .Y(n120) );
  OAI21X1 U122 ( .A(n121), .B(A[1]), .C(n154), .Y(n122) );
  NAND2X1 U123 ( .A(B[0]), .B(n153), .Y(n121) );
  OR2X2 U63 ( .A(A[31]), .B(B[30]), .Y(n63) );
  INVX2 U1 ( .A(n61), .Y(n123) );
  INVX2 U2 ( .A(A[15]), .Y(n124) );
  INVX2 U3 ( .A(A[16]), .Y(n125) );
  INVX2 U4 ( .A(A[17]), .Y(n126) );
  INVX2 U5 ( .A(A[18]), .Y(n127) );
  INVX2 U6 ( .A(A[19]), .Y(n128) );
  INVX2 U7 ( .A(A[20]), .Y(n129) );
  INVX2 U8 ( .A(A[21]), .Y(n130) );
  INVX2 U9 ( .A(A[22]), .Y(n131) );
  INVX2 U10 ( .A(A[23]), .Y(n132) );
  INVX2 U11 ( .A(A[24]), .Y(n133) );
  INVX2 U12 ( .A(A[25]), .Y(n134) );
  INVX2 U13 ( .A(A[26]), .Y(n135) );
  INVX2 U14 ( .A(A[27]), .Y(n136) );
  INVX2 U15 ( .A(A[28]), .Y(n137) );
  INVX2 U16 ( .A(A[29]), .Y(n138) );
  INVX2 U17 ( .A(A[31]), .Y(n139) );
  INVX2 U18 ( .A(A[14]), .Y(n140) );
  INVX2 U19 ( .A(A[13]), .Y(n141) );
  INVX2 U20 ( .A(A[12]), .Y(n142) );
  INVX2 U21 ( .A(A[11]), .Y(n143) );
  INVX2 U22 ( .A(A[9]), .Y(n144) );
  INVX2 U23 ( .A(A[8]), .Y(n145) );
  INVX2 U24 ( .A(A[7]), .Y(n146) );
  INVX2 U25 ( .A(A[6]), .Y(n147) );
  INVX2 U26 ( .A(A[5]), .Y(n148) );
  INVX2 U27 ( .A(A[4]), .Y(n149) );
  INVX2 U28 ( .A(A[3]), .Y(n150) );
  INVX2 U29 ( .A(A[2]), .Y(n151) );
  INVX2 U30 ( .A(n122), .Y(n152) );
  INVX2 U31 ( .A(A[0]), .Y(n153) );
  INVX2 U32 ( .A(B[1]), .Y(n154) );
  INVX2 U33 ( .A(B[2]), .Y(n155) );
  INVX2 U34 ( .A(B[3]), .Y(n156) );
  INVX2 U35 ( .A(B[4]), .Y(n157) );
  INVX2 U36 ( .A(B[5]), .Y(n158) );
  INVX2 U37 ( .A(B[6]), .Y(n159) );
  INVX2 U38 ( .A(B[7]), .Y(n160) );
  INVX2 U39 ( .A(B[8]), .Y(n161) );
  INVX2 U40 ( .A(B[10]), .Y(n162) );
  INVX2 U41 ( .A(B[11]), .Y(n163) );
  INVX2 U42 ( .A(B[12]), .Y(n164) );
  INVX2 U43 ( .A(B[13]), .Y(n165) );
  INVX2 U44 ( .A(B[14]), .Y(n166) );
  INVX2 U45 ( .A(B[15]), .Y(n167) );
  INVX2 U46 ( .A(B[16]), .Y(n168) );
  INVX2 U47 ( .A(B[17]), .Y(n169) );
  INVX2 U48 ( .A(B[18]), .Y(n170) );
  INVX2 U49 ( .A(B[19]), .Y(n171) );
  INVX2 U50 ( .A(B[20]), .Y(n172) );
  INVX2 U51 ( .A(B[21]), .Y(n173) );
  INVX2 U52 ( .A(B[22]), .Y(n174) );
  INVX2 U53 ( .A(B[23]), .Y(n175) );
  INVX2 U54 ( .A(B[24]), .Y(n176) );
  INVX2 U55 ( .A(B[25]), .Y(n177) );
  INVX2 U56 ( .A(B[26]), .Y(n178) );
  INVX2 U57 ( .A(B[27]), .Y(n179) );
  INVX2 U58 ( .A(B[28]), .Y(n180) );
  INVX2 U59 ( .A(B[29]), .Y(n181) );
  INVX2 U60 ( .A(B[31]), .Y(n182) );
endmodule


module CannyEdge_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n13), .B(\SUMB[5][5] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n53), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n23), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n31), .B(\SUMB[4][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n28), .B(\SUMB[4][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n29), .B(\SUMB[4][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n26), .B(\SUMB[6][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][2] ), .Y(n11) );
  AND2X2 U11 ( .A(n25), .B(\SUMB[6][3] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[4][5] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[7][4] ), .B(n10), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n9), .B(\SUMB[5][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n21), .B(\SUMB[3][1] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n15), .B(\SUMB[3][2] ), .Y(n31) );
  AND2X2 U31 ( .A(n20), .B(\ab[3][7] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n12), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n11), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n32), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n11), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n12), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n10), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n21), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n27), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n31), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n29), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n6), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n7), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n8), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n9), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n13), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n23), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n24), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n25), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n26), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n32), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n14), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n14), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n22), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n22), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n21), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n20), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n18), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n17), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n16), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n34), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n35), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n37), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n38), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n39), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n33), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n34), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n35), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n36), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n37), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n38), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n39), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n33), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n35), .B(\SUMB[6][4] ), .Y(n3) );
  AND2X2 U3 ( .A(n32), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n36), .B(\SUMB[2][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n37), .B(\SUMB[2][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[2][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n39), .B(\SUMB[2][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n40), .B(\SUMB[2][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n41), .B(\SUMB[2][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n27), .B(\SUMB[4][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n33), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n11), .B(n44), .Y(n14) );
  AND2X2 U14 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n21) );
  AND2X2 U21 ( .A(n4), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[3][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][5] ), .Y(n27) );
  AND2X2 U27 ( .A(n23), .B(\SUMB[4][1] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][2] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][3] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][4] ), .Y(n31) );
  AND2X2 U31 ( .A(n28), .B(\SUMB[5][1] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][2] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][3] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][4] ), .Y(n35) );
  AND2X2 U35 ( .A(n20), .B(\SUMB[1][1] ), .Y(n36) );
  AND2X2 U36 ( .A(n15), .B(\SUMB[1][2] ), .Y(n37) );
  AND2X2 U37 ( .A(n21), .B(\SUMB[1][3] ), .Y(n38) );
  AND2X2 U38 ( .A(n16), .B(\SUMB[1][4] ), .Y(n39) );
  AND2X2 U39 ( .A(n17), .B(\SUMB[1][5] ), .Y(n40) );
  AND2X2 U40 ( .A(n18), .B(\SUMB[1][6] ), .Y(n41) );
  AND2X2 U41 ( .A(n19), .B(\ab[1][7] ), .Y(n42) );
  XNOR2X1 U42 ( .A(n61), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U43 ( .A(n10), .B(n42), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][3] ), .B(n13), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][2] ), .B(n12), .Y(n46) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n14), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n14), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n20), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n15), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n21), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n16), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n17), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n18), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n19), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n36), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n37), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n38), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n39), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n40), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n41), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n5), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n6), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n7), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n8), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n9), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n42), .B(n10), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n23), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n24), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n25), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n26), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n27), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n28), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n29), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n30), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n31), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n44), .B(n11), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n32), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n33), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n34), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n35), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n46), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n46), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n45), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n45), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n22), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_4 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n12), .B(\SUMB[5][5] ), .Y(n3) );
  AND2X2 U3 ( .A(n22), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n26), .B(\SUMB[4][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n25), .B(\SUMB[6][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n23), .B(\SUMB[6][2] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][3] ), .Y(n11) );
  AND2X2 U11 ( .A(n30), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(\SUMB[7][4] ), .B(n9), .Y(n13) );
  AND2X2 U13 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(n4), .B(\SUMB[7][1] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[5][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][2] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][3] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][4] ), .Y(n25) );
  AND2X2 U25 ( .A(n14), .B(\SUMB[3][1] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n20), .B(\ab[3][7] ), .Y(n31) );
  XNOR2X1 U31 ( .A(n55), .B(n21), .Y(PRODUCT[9]) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n11), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n10), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n31), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n10), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n11), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n9), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n14), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n26), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n27), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n29), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n5), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n6), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n7), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n8), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n22), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n23), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n24), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n25), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n31), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n13), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n13), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n52), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n53), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n54), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n21), .Y(n36) );
  INVX2 U83 ( .A(n40), .Y(n52) );
  INVX2 U84 ( .A(n44), .Y(n53) );
  INVX2 U85 ( .A(n41), .Y(n54) );
  INVX2 U86 ( .A(\A1[7] ), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_6 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n12), .B(\SUMB[5][5] ), .Y(n3) );
  AND2X2 U3 ( .A(n22), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n26), .B(\SUMB[4][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n25), .B(\SUMB[6][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n23), .B(\SUMB[6][2] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][3] ), .Y(n11) );
  AND2X2 U11 ( .A(n30), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(\SUMB[7][4] ), .B(n9), .Y(n13) );
  AND2X2 U13 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(n4), .B(\SUMB[7][1] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[5][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][2] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][3] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][4] ), .Y(n25) );
  AND2X2 U25 ( .A(n14), .B(\SUMB[3][1] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n20), .B(\ab[3][7] ), .Y(n31) );
  XNOR2X1 U31 ( .A(n53), .B(n21), .Y(PRODUCT[9]) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n11), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n10), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n31), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n10), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n11), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n9), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n14), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n26), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n27), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n29), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n5), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n6), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n7), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n8), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n22), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n23), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n24), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n25), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n31), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n13), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n13), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n21), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_8 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n36), .B(\SUMB[6][4] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n33), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n37), .B(\SUMB[2][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[2][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n39), .B(\SUMB[2][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n40), .B(\SUMB[2][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n41), .B(\SUMB[2][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n42), .B(\SUMB[2][6] ), .Y(n11) );
  AND2X2 U11 ( .A(n28), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n35), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(n12), .B(n44), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[3][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[4][4] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][1] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][2] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][3] ), .Y(n35) );
  AND2X2 U35 ( .A(n32), .B(\SUMB[5][4] ), .Y(n36) );
  AND2X2 U36 ( .A(n22), .B(\SUMB[1][1] ), .Y(n37) );
  AND2X2 U37 ( .A(n16), .B(\SUMB[1][2] ), .Y(n38) );
  AND2X2 U38 ( .A(n17), .B(\SUMB[1][3] ), .Y(n39) );
  AND2X2 U39 ( .A(n18), .B(\SUMB[1][4] ), .Y(n40) );
  AND2X2 U40 ( .A(n19), .B(\SUMB[1][5] ), .Y(n41) );
  AND2X2 U41 ( .A(n20), .B(\SUMB[1][6] ), .Y(n42) );
  AND2X2 U42 ( .A(n21), .B(\ab[1][7] ), .Y(n43) );
  AND2X2 U43 ( .A(n11), .B(n43), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][3] ), .B(n14), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][2] ), .B(n13), .Y(n46) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n15), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n15), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n22), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n16), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n17), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n18), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n19), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n20), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n21), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n37), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n38), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n39), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n40), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n41), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n42), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n6), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n7), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n8), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n9), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n10), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n43), .B(n11), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n24), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n25), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n26), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n27), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n28), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n29), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n30), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n31), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n32), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n44), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n33), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n34), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n35), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n36), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n46), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n46), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n45), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n45), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n23), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_9 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n22), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n21), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n20), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n19), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n18), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n17), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n34), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n35), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n37), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n38), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n39), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n33), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n34), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n35), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n36), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n37), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n38), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n39), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n33), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW02_mult_10 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n13), .B(\SUMB[5][5] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n53), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n23), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n30), .B(\SUMB[4][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n26), .B(\SUMB[6][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][2] ), .Y(n11) );
  AND2X2 U11 ( .A(n25), .B(\SUMB[6][3] ), .Y(n12) );
  AND2X2 U12 ( .A(n31), .B(\SUMB[4][5] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[7][4] ), .B(n10), .Y(n14) );
  AND2X2 U14 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n15) );
  AND2X2 U15 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n20) );
  AND2X2 U20 ( .A(n20), .B(\ab[3][6] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n9), .B(\SUMB[5][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][1] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][2] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][4] ), .Y(n30) );
  AND2X2 U30 ( .A(n19), .B(\SUMB[3][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n21), .B(\ab[3][7] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n12), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n11), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n32), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n11), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n12), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n10), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n15), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n16), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n17), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n18), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n19), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n20), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n27), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n28), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n29), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n30), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n31), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n21), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n6), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n7), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n8), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n9), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n13), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n23), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n24), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n25), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n26), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n32), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n14), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n14), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n22), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_11 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [7:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , n3, n4, n5, n6, n7, n8, n9, n22, n20, n18, n16, n14,
         n12, n10, \ab[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[30][1] ,
         \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] ,
         \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[30][0] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] ,
         \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][5] , \CARRYB[25][4] ,
         \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] ,
         \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] ,
         \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][6] ,
         \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] ,
         \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] ,
         \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][6] ,
         \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] ,
         \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] ,
         \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \CARRYB[15][6] ,
         \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] ,
         \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][6] ,
         \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] ,
         \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50;

  AND2X2 U2 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n3) );
  AND2X2 U3 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n4) );
  AND2X2 U4 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n5) );
  AND2X2 U5 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n6) );
  AND2X2 U6 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n7) );
  AND2X2 U7 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n8) );
  AND2X2 U8 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n9) );
  XOR2X1 U24 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U25 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U26 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U27 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U28 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U29 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U30 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  NOR2X1 U41 ( .A(n50), .B(n42), .Y(\ab[1][7] ) );
  NOR2X1 U42 ( .A(n49), .B(n42), .Y(\ab[1][6] ) );
  NOR2X1 U43 ( .A(n48), .B(n42), .Y(\ab[1][5] ) );
  NOR2X1 U44 ( .A(n47), .B(n42), .Y(\ab[1][4] ) );
  NOR2X1 U45 ( .A(n46), .B(n42), .Y(\ab[1][3] ) );
  NOR2X1 U46 ( .A(n45), .B(n42), .Y(\ab[1][2] ) );
  NOR2X1 U47 ( .A(n44), .B(n42), .Y(\ab[1][1] ) );
  NOR2X1 U48 ( .A(n43), .B(n42), .Y(\ab[1][0] ) );
  NOR2X1 U49 ( .A(n50), .B(n41), .Y(\ab[0][7] ) );
  NOR2X1 U50 ( .A(n49), .B(n41), .Y(\ab[0][6] ) );
  NOR2X1 U51 ( .A(n48), .B(n41), .Y(\ab[0][5] ) );
  NOR2X1 U52 ( .A(n47), .B(n41), .Y(\ab[0][4] ) );
  NOR2X1 U53 ( .A(n46), .B(n41), .Y(\ab[0][3] ) );
  NOR2X1 U54 ( .A(n45), .B(n41), .Y(\ab[0][2] ) );
  NOR2X1 U55 ( .A(n44), .B(n41), .Y(\ab[0][1] ) );
  NOR2X1 U56 ( .A(n43), .B(n41), .Y(PRODUCT[0]) );
  FAX1 S4_0 ( .A(n34), .B(\CARRYB[30][0] ), .C(\SUMB[30][1] ), .YS(PRODUCT[31]) );
  FAX1 S1_30_0 ( .A(n34), .B(\CARRYB[29][0] ), .C(\SUMB[29][1] ), .YC(
        \CARRYB[30][0] ), .YS(PRODUCT[30]) );
  FAX1 S1_29_0 ( .A(n34), .B(\CARRYB[28][0] ), .C(\SUMB[28][1] ), .YC(
        \CARRYB[29][0] ), .YS(PRODUCT[29]) );
  FAX1 S1_28_0 ( .A(n34), .B(\CARRYB[27][0] ), .C(\SUMB[27][1] ), .YC(
        \CARRYB[28][0] ), .YS(PRODUCT[28]) );
  FAX1 S1_27_0 ( .A(n34), .B(\CARRYB[26][0] ), .C(\SUMB[26][1] ), .YC(
        \CARRYB[27][0] ), .YS(PRODUCT[27]) );
  FAX1 S1_26_0 ( .A(n34), .B(\CARRYB[25][0] ), .C(\SUMB[25][1] ), .YC(
        \CARRYB[26][0] ), .YS(PRODUCT[26]) );
  FAX1 S1_25_0 ( .A(n34), .B(\CARRYB[24][0] ), .C(\SUMB[24][1] ), .YC(
        \CARRYB[25][0] ), .YS(PRODUCT[25]) );
  FAX1 S1_24_0 ( .A(n34), .B(\CARRYB[23][0] ), .C(\SUMB[23][1] ), .YC(
        \CARRYB[24][0] ), .YS(PRODUCT[24]) );
  FAX1 S1_23_0 ( .A(n34), .B(\CARRYB[22][0] ), .C(\SUMB[22][1] ), .YC(
        \CARRYB[23][0] ), .YS(PRODUCT[23]) );
  FAX1 S1_22_0 ( .A(n34), .B(\CARRYB[21][0] ), .C(\SUMB[21][1] ), .YC(
        \CARRYB[22][0] ), .YS(PRODUCT[22]) );
  FAX1 S1_21_0 ( .A(n34), .B(\CARRYB[20][0] ), .C(\SUMB[20][1] ), .YC(
        \CARRYB[21][0] ), .YS(PRODUCT[21]) );
  FAX1 S1_20_0 ( .A(n34), .B(\CARRYB[19][0] ), .C(\SUMB[19][1] ), .YC(
        \CARRYB[20][0] ), .YS(PRODUCT[20]) );
  FAX1 S1_19_0 ( .A(n34), .B(\CARRYB[18][0] ), .C(\SUMB[18][1] ), .YC(
        \CARRYB[19][0] ), .YS(PRODUCT[19]) );
  FAX1 S1_18_0 ( .A(n34), .B(\CARRYB[17][0] ), .C(\SUMB[17][1] ), .YC(
        \CARRYB[18][0] ), .YS(PRODUCT[18]) );
  FAX1 S1_17_0 ( .A(n34), .B(\CARRYB[16][0] ), .C(\SUMB[16][1] ), .YC(
        \CARRYB[17][0] ), .YS(PRODUCT[17]) );
  FAX1 S1_16_0 ( .A(n34), .B(\CARRYB[15][0] ), .C(\SUMB[15][1] ), .YC(
        \CARRYB[16][0] ), .YS(PRODUCT[16]) );
  FAX1 S1_15_0 ( .A(n34), .B(\CARRYB[14][0] ), .C(\SUMB[14][1] ), .YC(
        \CARRYB[15][0] ), .YS(PRODUCT[15]) );
  FAX1 S1_14_0 ( .A(n34), .B(\CARRYB[13][0] ), .C(\SUMB[13][1] ), .YC(
        \CARRYB[14][0] ), .YS(PRODUCT[14]) );
  FAX1 S1_13_0 ( .A(n34), .B(\CARRYB[12][0] ), .C(\SUMB[12][1] ), .YC(
        \CARRYB[13][0] ), .YS(PRODUCT[13]) );
  FAX1 S1_12_0 ( .A(n34), .B(\CARRYB[11][0] ), .C(\SUMB[11][1] ), .YC(
        \CARRYB[12][0] ), .YS(PRODUCT[12]) );
  FAX1 S1_11_0 ( .A(n34), .B(\CARRYB[10][0] ), .C(\SUMB[10][1] ), .YC(
        \CARRYB[11][0] ), .YS(PRODUCT[11]) );
  FAX1 S1_10_0 ( .A(n34), .B(\CARRYB[9][0] ), .C(\SUMB[9][1] ), .YC(
        \CARRYB[10][0] ), .YS(PRODUCT[10]) );
  FAX1 S1_9_0 ( .A(n34), .B(\CARRYB[8][0] ), .C(\SUMB[8][1] ), .YC(
        \CARRYB[9][0] ), .YS(PRODUCT[9]) );
  FAX1 S1_8_0 ( .A(n34), .B(\CARRYB[7][0] ), .C(\SUMB[7][1] ), .YC(
        \CARRYB[8][0] ), .YS(PRODUCT[8]) );
  FAX1 S1_7_0 ( .A(n34), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(PRODUCT[7]) );
  FAX1 S1_6_0 ( .A(n34), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(PRODUCT[6]) );
  FAX1 S1_5_0 ( .A(n34), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(PRODUCT[5]) );
  FAX1 S1_4_0 ( .A(n34), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(PRODUCT[4]) );
  FAX1 S1_3_0 ( .A(n34), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(PRODUCT[3]) );
  FAX1 S1_2_0 ( .A(n34), .B(n9), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), .YS(
        PRODUCT[2]) );
  NAND2X1 U22 ( .A(B[0]), .B(A[9]), .Y(n22) );
  FAX1 S2_30_1 ( .A(n36), .B(\CARRYB[29][1] ), .C(\SUMB[29][2] ), .YS(
        \SUMB[30][1] ) );
  FAX1 S2_29_1 ( .A(n36), .B(\CARRYB[28][1] ), .C(\SUMB[28][2] ), .YC(
        \CARRYB[29][1] ), .YS(\SUMB[29][1] ) );
  FAX1 S2_28_1 ( .A(n36), .B(\CARRYB[27][1] ), .C(\SUMB[27][2] ), .YC(
        \CARRYB[28][1] ), .YS(\SUMB[28][1] ) );
  FAX1 S2_27_1 ( .A(n36), .B(\CARRYB[26][1] ), .C(\SUMB[26][2] ), .YC(
        \CARRYB[27][1] ), .YS(\SUMB[27][1] ) );
  FAX1 S2_26_1 ( .A(n36), .B(\CARRYB[25][1] ), .C(\SUMB[25][2] ), .YC(
        \CARRYB[26][1] ), .YS(\SUMB[26][1] ) );
  FAX1 S2_25_1 ( .A(n36), .B(\CARRYB[24][1] ), .C(\SUMB[24][2] ), .YC(
        \CARRYB[25][1] ), .YS(\SUMB[25][1] ) );
  FAX1 S2_24_1 ( .A(n36), .B(\CARRYB[23][1] ), .C(\SUMB[23][2] ), .YC(
        \CARRYB[24][1] ), .YS(\SUMB[24][1] ) );
  FAX1 S2_23_1 ( .A(n36), .B(\CARRYB[22][1] ), .C(\SUMB[22][2] ), .YC(
        \CARRYB[23][1] ), .YS(\SUMB[23][1] ) );
  FAX1 S2_22_1 ( .A(n36), .B(\CARRYB[21][1] ), .C(\SUMB[21][2] ), .YC(
        \CARRYB[22][1] ), .YS(\SUMB[22][1] ) );
  FAX1 S2_21_1 ( .A(n36), .B(\CARRYB[20][1] ), .C(\SUMB[20][2] ), .YC(
        \CARRYB[21][1] ), .YS(\SUMB[21][1] ) );
  FAX1 S2_20_1 ( .A(n36), .B(\CARRYB[19][1] ), .C(\SUMB[19][2] ), .YC(
        \CARRYB[20][1] ), .YS(\SUMB[20][1] ) );
  FAX1 S2_19_1 ( .A(n36), .B(\CARRYB[18][1] ), .C(\SUMB[18][2] ), .YC(
        \CARRYB[19][1] ), .YS(\SUMB[19][1] ) );
  FAX1 S2_18_1 ( .A(n36), .B(\CARRYB[17][1] ), .C(\SUMB[17][2] ), .YC(
        \CARRYB[18][1] ), .YS(\SUMB[18][1] ) );
  FAX1 S2_17_1 ( .A(n36), .B(\CARRYB[16][1] ), .C(\SUMB[16][2] ), .YC(
        \CARRYB[17][1] ), .YS(\SUMB[17][1] ) );
  FAX1 S2_16_1 ( .A(n36), .B(\CARRYB[15][1] ), .C(\SUMB[15][2] ), .YC(
        \CARRYB[16][1] ), .YS(\SUMB[16][1] ) );
  FAX1 S2_15_1 ( .A(n36), .B(\CARRYB[14][1] ), .C(\SUMB[14][2] ), .YC(
        \CARRYB[15][1] ), .YS(\SUMB[15][1] ) );
  FAX1 S2_14_1 ( .A(n36), .B(\CARRYB[13][1] ), .C(\SUMB[13][2] ), .YC(
        \CARRYB[14][1] ), .YS(\SUMB[14][1] ) );
  FAX1 S2_13_1 ( .A(n36), .B(\CARRYB[12][1] ), .C(\SUMB[12][2] ), .YC(
        \CARRYB[13][1] ), .YS(\SUMB[13][1] ) );
  FAX1 S2_12_1 ( .A(n36), .B(\CARRYB[11][1] ), .C(\SUMB[11][2] ), .YC(
        \CARRYB[12][1] ), .YS(\SUMB[12][1] ) );
  FAX1 S2_11_1 ( .A(n36), .B(\CARRYB[10][1] ), .C(\SUMB[10][2] ), .YC(
        \CARRYB[11][1] ), .YS(\SUMB[11][1] ) );
  FAX1 S2_10_1 ( .A(n36), .B(\CARRYB[9][1] ), .C(\SUMB[9][2] ), .YC(
        \CARRYB[10][1] ), .YS(\SUMB[10][1] ) );
  FAX1 S2_9_1 ( .A(n36), .B(\CARRYB[8][1] ), .C(\SUMB[8][2] ), .YC(
        \CARRYB[9][1] ), .YS(\SUMB[9][1] ) );
  FAX1 S2_8_1 ( .A(n36), .B(\CARRYB[7][1] ), .C(\SUMB[7][2] ), .YC(
        \CARRYB[8][1] ), .YS(\SUMB[8][1] ) );
  FAX1 S2_7_1 ( .A(n36), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S2_6_1 ( .A(n36), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_5_1 ( .A(n36), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_4_1 ( .A(n36), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_3_1 ( .A(n36), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_2_1 ( .A(n36), .B(n8), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), .YS(
        \SUMB[2][1] ) );
  NAND2X1 U18 ( .A(B[1]), .B(A[9]), .Y(n18) );
  FAX1 S2_29_2 ( .A(n38), .B(\CARRYB[28][2] ), .C(\SUMB[28][3] ), .YS(
        \SUMB[29][2] ) );
  FAX1 S2_28_2 ( .A(n38), .B(\CARRYB[27][2] ), .C(\SUMB[27][3] ), .YC(
        \CARRYB[28][2] ), .YS(\SUMB[28][2] ) );
  FAX1 S2_27_2 ( .A(n38), .B(\CARRYB[26][2] ), .C(\SUMB[26][3] ), .YC(
        \CARRYB[27][2] ), .YS(\SUMB[27][2] ) );
  FAX1 S2_26_2 ( .A(n38), .B(\CARRYB[25][2] ), .C(\SUMB[25][3] ), .YC(
        \CARRYB[26][2] ), .YS(\SUMB[26][2] ) );
  FAX1 S2_25_2 ( .A(n38), .B(\CARRYB[24][2] ), .C(\SUMB[24][3] ), .YC(
        \CARRYB[25][2] ), .YS(\SUMB[25][2] ) );
  FAX1 S2_24_2 ( .A(n38), .B(\CARRYB[23][2] ), .C(\SUMB[23][3] ), .YC(
        \CARRYB[24][2] ), .YS(\SUMB[24][2] ) );
  FAX1 S2_23_2 ( .A(n38), .B(\CARRYB[22][2] ), .C(\SUMB[22][3] ), .YC(
        \CARRYB[23][2] ), .YS(\SUMB[23][2] ) );
  FAX1 S2_22_2 ( .A(n38), .B(\CARRYB[21][2] ), .C(\SUMB[21][3] ), .YC(
        \CARRYB[22][2] ), .YS(\SUMB[22][2] ) );
  FAX1 S2_21_2 ( .A(n38), .B(\CARRYB[20][2] ), .C(\SUMB[20][3] ), .YC(
        \CARRYB[21][2] ), .YS(\SUMB[21][2] ) );
  FAX1 S2_20_2 ( .A(n38), .B(\CARRYB[19][2] ), .C(\SUMB[19][3] ), .YC(
        \CARRYB[20][2] ), .YS(\SUMB[20][2] ) );
  FAX1 S2_19_2 ( .A(n38), .B(\CARRYB[18][2] ), .C(\SUMB[18][3] ), .YC(
        \CARRYB[19][2] ), .YS(\SUMB[19][2] ) );
  FAX1 S2_18_2 ( .A(n38), .B(\CARRYB[17][2] ), .C(\SUMB[17][3] ), .YC(
        \CARRYB[18][2] ), .YS(\SUMB[18][2] ) );
  FAX1 S2_17_2 ( .A(n38), .B(\CARRYB[16][2] ), .C(\SUMB[16][3] ), .YC(
        \CARRYB[17][2] ), .YS(\SUMB[17][2] ) );
  FAX1 S2_16_2 ( .A(n38), .B(\CARRYB[15][2] ), .C(\SUMB[15][3] ), .YC(
        \CARRYB[16][2] ), .YS(\SUMB[16][2] ) );
  FAX1 S2_15_2 ( .A(n38), .B(\CARRYB[14][2] ), .C(\SUMB[14][3] ), .YC(
        \CARRYB[15][2] ), .YS(\SUMB[15][2] ) );
  FAX1 S2_14_2 ( .A(n38), .B(\CARRYB[13][2] ), .C(\SUMB[13][3] ), .YC(
        \CARRYB[14][2] ), .YS(\SUMB[14][2] ) );
  FAX1 S2_13_2 ( .A(n38), .B(\CARRYB[12][2] ), .C(\SUMB[12][3] ), .YC(
        \CARRYB[13][2] ), .YS(\SUMB[13][2] ) );
  FAX1 S2_12_2 ( .A(n38), .B(\CARRYB[11][2] ), .C(\SUMB[11][3] ), .YC(
        \CARRYB[12][2] ), .YS(\SUMB[12][2] ) );
  FAX1 S2_11_2 ( .A(n38), .B(\CARRYB[10][2] ), .C(\SUMB[10][3] ), .YC(
        \CARRYB[11][2] ), .YS(\SUMB[11][2] ) );
  FAX1 S2_10_2 ( .A(n38), .B(\CARRYB[9][2] ), .C(\SUMB[9][3] ), .YC(
        \CARRYB[10][2] ), .YS(\SUMB[10][2] ) );
  FAX1 S2_9_2 ( .A(n38), .B(\CARRYB[8][2] ), .C(\SUMB[8][3] ), .YC(
        \CARRYB[9][2] ), .YS(\SUMB[9][2] ) );
  FAX1 S2_8_2 ( .A(n38), .B(\CARRYB[7][2] ), .C(\SUMB[7][3] ), .YC(
        \CARRYB[8][2] ), .YS(\SUMB[8][2] ) );
  FAX1 S2_7_2 ( .A(n38), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(n38), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_5_2 ( .A(n38), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_4_2 ( .A(n38), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_3_2 ( .A(n38), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_2_2 ( .A(n38), .B(n7), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), .YS(
        \SUMB[2][2] ) );
  NAND2X1 U14 ( .A(B[2]), .B(A[9]), .Y(n14) );
  FAX1 S2_28_3 ( .A(n35), .B(\CARRYB[27][3] ), .C(\SUMB[27][4] ), .YS(
        \SUMB[28][3] ) );
  FAX1 S2_27_3 ( .A(n35), .B(\CARRYB[26][3] ), .C(\SUMB[26][4] ), .YC(
        \CARRYB[27][3] ), .YS(\SUMB[27][3] ) );
  FAX1 S2_26_3 ( .A(n35), .B(\CARRYB[25][3] ), .C(\SUMB[25][4] ), .YC(
        \CARRYB[26][3] ), .YS(\SUMB[26][3] ) );
  FAX1 S2_25_3 ( .A(n35), .B(\CARRYB[24][3] ), .C(\SUMB[24][4] ), .YC(
        \CARRYB[25][3] ), .YS(\SUMB[25][3] ) );
  FAX1 S2_24_3 ( .A(n35), .B(\CARRYB[23][3] ), .C(\SUMB[23][4] ), .YC(
        \CARRYB[24][3] ), .YS(\SUMB[24][3] ) );
  FAX1 S2_23_3 ( .A(n35), .B(\CARRYB[22][3] ), .C(\SUMB[22][4] ), .YC(
        \CARRYB[23][3] ), .YS(\SUMB[23][3] ) );
  FAX1 S2_22_3 ( .A(n35), .B(\CARRYB[21][3] ), .C(\SUMB[21][4] ), .YC(
        \CARRYB[22][3] ), .YS(\SUMB[22][3] ) );
  FAX1 S2_21_3 ( .A(n35), .B(\CARRYB[20][3] ), .C(\SUMB[20][4] ), .YC(
        \CARRYB[21][3] ), .YS(\SUMB[21][3] ) );
  FAX1 S2_20_3 ( .A(n35), .B(\CARRYB[19][3] ), .C(\SUMB[19][4] ), .YC(
        \CARRYB[20][3] ), .YS(\SUMB[20][3] ) );
  FAX1 S2_19_3 ( .A(n35), .B(\CARRYB[18][3] ), .C(\SUMB[18][4] ), .YC(
        \CARRYB[19][3] ), .YS(\SUMB[19][3] ) );
  FAX1 S2_18_3 ( .A(n35), .B(\CARRYB[17][3] ), .C(\SUMB[17][4] ), .YC(
        \CARRYB[18][3] ), .YS(\SUMB[18][3] ) );
  FAX1 S2_17_3 ( .A(n35), .B(\CARRYB[16][3] ), .C(\SUMB[16][4] ), .YC(
        \CARRYB[17][3] ), .YS(\SUMB[17][3] ) );
  FAX1 S2_16_3 ( .A(n35), .B(\CARRYB[15][3] ), .C(\SUMB[15][4] ), .YC(
        \CARRYB[16][3] ), .YS(\SUMB[16][3] ) );
  FAX1 S2_15_3 ( .A(n35), .B(\CARRYB[14][3] ), .C(\SUMB[14][4] ), .YC(
        \CARRYB[15][3] ), .YS(\SUMB[15][3] ) );
  FAX1 S2_14_3 ( .A(n35), .B(\CARRYB[13][3] ), .C(\SUMB[13][4] ), .YC(
        \CARRYB[14][3] ), .YS(\SUMB[14][3] ) );
  FAX1 S2_13_3 ( .A(n35), .B(\CARRYB[12][3] ), .C(\SUMB[12][4] ), .YC(
        \CARRYB[13][3] ), .YS(\SUMB[13][3] ) );
  FAX1 S2_12_3 ( .A(n35), .B(\CARRYB[11][3] ), .C(\SUMB[11][4] ), .YC(
        \CARRYB[12][3] ), .YS(\SUMB[12][3] ) );
  FAX1 S2_11_3 ( .A(n35), .B(\CARRYB[10][3] ), .C(\SUMB[10][4] ), .YC(
        \CARRYB[11][3] ), .YS(\SUMB[11][3] ) );
  FAX1 S2_10_3 ( .A(n35), .B(\CARRYB[9][3] ), .C(\SUMB[9][4] ), .YC(
        \CARRYB[10][3] ), .YS(\SUMB[10][3] ) );
  FAX1 S2_9_3 ( .A(n35), .B(\CARRYB[8][3] ), .C(\SUMB[8][4] ), .YC(
        \CARRYB[9][3] ), .YS(\SUMB[9][3] ) );
  FAX1 S2_8_3 ( .A(n35), .B(\CARRYB[7][3] ), .C(\SUMB[7][4] ), .YC(
        \CARRYB[8][3] ), .YS(\SUMB[8][3] ) );
  FAX1 S2_7_3 ( .A(n35), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(n35), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(n35), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_4_3 ( .A(n35), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_3_3 ( .A(n35), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_2_3 ( .A(n35), .B(n6), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), .YS(
        \SUMB[2][3] ) );
  NAND2X1 U20 ( .A(B[3]), .B(A[9]), .Y(n20) );
  FAX1 S2_27_4 ( .A(n37), .B(\CARRYB[26][4] ), .C(\SUMB[26][5] ), .YS(
        \SUMB[27][4] ) );
  FAX1 S2_26_4 ( .A(n37), .B(\CARRYB[25][4] ), .C(\SUMB[25][5] ), .YC(
        \CARRYB[26][4] ), .YS(\SUMB[26][4] ) );
  FAX1 S2_25_4 ( .A(n37), .B(\CARRYB[24][4] ), .C(\SUMB[24][5] ), .YC(
        \CARRYB[25][4] ), .YS(\SUMB[25][4] ) );
  FAX1 S2_24_4 ( .A(n37), .B(\CARRYB[23][4] ), .C(\SUMB[23][5] ), .YC(
        \CARRYB[24][4] ), .YS(\SUMB[24][4] ) );
  FAX1 S2_23_4 ( .A(n37), .B(\CARRYB[22][4] ), .C(\SUMB[22][5] ), .YC(
        \CARRYB[23][4] ), .YS(\SUMB[23][4] ) );
  FAX1 S2_22_4 ( .A(n37), .B(\CARRYB[21][4] ), .C(\SUMB[21][5] ), .YC(
        \CARRYB[22][4] ), .YS(\SUMB[22][4] ) );
  FAX1 S2_21_4 ( .A(n37), .B(\CARRYB[20][4] ), .C(\SUMB[20][5] ), .YC(
        \CARRYB[21][4] ), .YS(\SUMB[21][4] ) );
  FAX1 S2_20_4 ( .A(n37), .B(\CARRYB[19][4] ), .C(\SUMB[19][5] ), .YC(
        \CARRYB[20][4] ), .YS(\SUMB[20][4] ) );
  FAX1 S2_19_4 ( .A(n37), .B(\CARRYB[18][4] ), .C(\SUMB[18][5] ), .YC(
        \CARRYB[19][4] ), .YS(\SUMB[19][4] ) );
  FAX1 S2_18_4 ( .A(n37), .B(\CARRYB[17][4] ), .C(\SUMB[17][5] ), .YC(
        \CARRYB[18][4] ), .YS(\SUMB[18][4] ) );
  FAX1 S2_17_4 ( .A(n37), .B(\CARRYB[16][4] ), .C(\SUMB[16][5] ), .YC(
        \CARRYB[17][4] ), .YS(\SUMB[17][4] ) );
  FAX1 S2_16_4 ( .A(n37), .B(\CARRYB[15][4] ), .C(\SUMB[15][5] ), .YC(
        \CARRYB[16][4] ), .YS(\SUMB[16][4] ) );
  FAX1 S2_15_4 ( .A(n37), .B(\CARRYB[14][4] ), .C(\SUMB[14][5] ), .YC(
        \CARRYB[15][4] ), .YS(\SUMB[15][4] ) );
  FAX1 S2_14_4 ( .A(n37), .B(\CARRYB[13][4] ), .C(\SUMB[13][5] ), .YC(
        \CARRYB[14][4] ), .YS(\SUMB[14][4] ) );
  FAX1 S2_13_4 ( .A(n37), .B(\CARRYB[12][4] ), .C(\SUMB[12][5] ), .YC(
        \CARRYB[13][4] ), .YS(\SUMB[13][4] ) );
  FAX1 S2_12_4 ( .A(n37), .B(\CARRYB[11][4] ), .C(\SUMB[11][5] ), .YC(
        \CARRYB[12][4] ), .YS(\SUMB[12][4] ) );
  FAX1 S2_11_4 ( .A(n37), .B(\CARRYB[10][4] ), .C(\SUMB[10][5] ), .YC(
        \CARRYB[11][4] ), .YS(\SUMB[11][4] ) );
  FAX1 S2_10_4 ( .A(n37), .B(\CARRYB[9][4] ), .C(\SUMB[9][5] ), .YC(
        \CARRYB[10][4] ), .YS(\SUMB[10][4] ) );
  FAX1 S2_9_4 ( .A(n37), .B(\CARRYB[8][4] ), .C(\SUMB[8][5] ), .YC(
        \CARRYB[9][4] ), .YS(\SUMB[9][4] ) );
  FAX1 S2_8_4 ( .A(n37), .B(\CARRYB[7][4] ), .C(\SUMB[7][5] ), .YC(
        \CARRYB[8][4] ), .YS(\SUMB[8][4] ) );
  FAX1 S2_7_4 ( .A(n37), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(n37), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(n37), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(n37), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_3_4 ( .A(n37), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_2_4 ( .A(n37), .B(n5), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), .YS(
        \SUMB[2][4] ) );
  NAND2X1 U16 ( .A(B[4]), .B(A[9]), .Y(n16) );
  FAX1 S2_26_5 ( .A(n39), .B(\CARRYB[25][5] ), .C(\SUMB[25][6] ), .YS(
        \SUMB[26][5] ) );
  FAX1 S3_25_6 ( .A(n40), .B(\CARRYB[24][6] ), .C(\ab[9][7] ), .YS(
        \SUMB[25][6] ) );
  FAX1 S2_25_5 ( .A(n39), .B(\CARRYB[24][5] ), .C(\SUMB[24][6] ), .YC(
        \CARRYB[25][5] ), .YS(\SUMB[25][5] ) );
  FAX1 S3_24_6 ( .A(n40), .B(\CARRYB[23][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[24][6] ), .YS(\SUMB[24][6] ) );
  FAX1 S2_24_5 ( .A(n39), .B(\CARRYB[23][5] ), .C(\SUMB[23][6] ), .YC(
        \CARRYB[24][5] ), .YS(\SUMB[24][5] ) );
  FAX1 S3_23_6 ( .A(n40), .B(\CARRYB[22][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[23][6] ), .YS(\SUMB[23][6] ) );
  FAX1 S2_23_5 ( .A(n39), .B(\CARRYB[22][5] ), .C(\SUMB[22][6] ), .YC(
        \CARRYB[23][5] ), .YS(\SUMB[23][5] ) );
  FAX1 S3_22_6 ( .A(n40), .B(\CARRYB[21][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[22][6] ), .YS(\SUMB[22][6] ) );
  FAX1 S2_22_5 ( .A(n39), .B(\CARRYB[21][5] ), .C(\SUMB[21][6] ), .YC(
        \CARRYB[22][5] ), .YS(\SUMB[22][5] ) );
  FAX1 S3_21_6 ( .A(n40), .B(\CARRYB[20][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[21][6] ), .YS(\SUMB[21][6] ) );
  FAX1 S2_21_5 ( .A(n39), .B(\CARRYB[20][5] ), .C(\SUMB[20][6] ), .YC(
        \CARRYB[21][5] ), .YS(\SUMB[21][5] ) );
  FAX1 S3_20_6 ( .A(n40), .B(\CARRYB[19][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[20][6] ), .YS(\SUMB[20][6] ) );
  FAX1 S2_20_5 ( .A(n39), .B(\CARRYB[19][5] ), .C(\SUMB[19][6] ), .YC(
        \CARRYB[20][5] ), .YS(\SUMB[20][5] ) );
  FAX1 S3_19_6 ( .A(n40), .B(\CARRYB[18][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[19][6] ), .YS(\SUMB[19][6] ) );
  FAX1 S2_19_5 ( .A(n39), .B(\CARRYB[18][5] ), .C(\SUMB[18][6] ), .YC(
        \CARRYB[19][5] ), .YS(\SUMB[19][5] ) );
  FAX1 S3_18_6 ( .A(n40), .B(\CARRYB[17][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[18][6] ), .YS(\SUMB[18][6] ) );
  FAX1 S2_18_5 ( .A(n39), .B(\CARRYB[17][5] ), .C(\SUMB[17][6] ), .YC(
        \CARRYB[18][5] ), .YS(\SUMB[18][5] ) );
  FAX1 S3_17_6 ( .A(n40), .B(\CARRYB[16][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[17][6] ), .YS(\SUMB[17][6] ) );
  FAX1 S2_17_5 ( .A(n39), .B(\CARRYB[16][5] ), .C(\SUMB[16][6] ), .YC(
        \CARRYB[17][5] ), .YS(\SUMB[17][5] ) );
  FAX1 S3_16_6 ( .A(n40), .B(\CARRYB[15][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[16][6] ), .YS(\SUMB[16][6] ) );
  FAX1 S2_16_5 ( .A(n39), .B(\CARRYB[15][5] ), .C(\SUMB[15][6] ), .YC(
        \CARRYB[16][5] ), .YS(\SUMB[16][5] ) );
  FAX1 S3_15_6 ( .A(n40), .B(\CARRYB[14][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[15][6] ), .YS(\SUMB[15][6] ) );
  FAX1 S2_15_5 ( .A(n39), .B(\CARRYB[14][5] ), .C(\SUMB[14][6] ), .YC(
        \CARRYB[15][5] ), .YS(\SUMB[15][5] ) );
  FAX1 S3_14_6 ( .A(n40), .B(\CARRYB[13][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[14][6] ), .YS(\SUMB[14][6] ) );
  FAX1 S2_14_5 ( .A(n39), .B(\CARRYB[13][5] ), .C(\SUMB[13][6] ), .YC(
        \CARRYB[14][5] ), .YS(\SUMB[14][5] ) );
  FAX1 S3_13_6 ( .A(n40), .B(\CARRYB[12][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[13][6] ), .YS(\SUMB[13][6] ) );
  FAX1 S2_13_5 ( .A(n39), .B(\CARRYB[12][5] ), .C(\SUMB[12][6] ), .YC(
        \CARRYB[13][5] ), .YS(\SUMB[13][5] ) );
  FAX1 S3_12_6 ( .A(n40), .B(\CARRYB[11][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[12][6] ), .YS(\SUMB[12][6] ) );
  FAX1 S2_12_5 ( .A(n39), .B(\CARRYB[11][5] ), .C(\SUMB[11][6] ), .YC(
        \CARRYB[12][5] ), .YS(\SUMB[12][5] ) );
  FAX1 S3_11_6 ( .A(n40), .B(\CARRYB[10][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[11][6] ), .YS(\SUMB[11][6] ) );
  FAX1 S2_11_5 ( .A(n39), .B(\CARRYB[10][5] ), .C(\SUMB[10][6] ), .YC(
        \CARRYB[11][5] ), .YS(\SUMB[11][5] ) );
  FAX1 S3_10_6 ( .A(n40), .B(\CARRYB[9][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[10][6] ), .YS(\SUMB[10][6] ) );
  FAX1 S2_10_5 ( .A(n39), .B(\CARRYB[9][5] ), .C(\SUMB[9][6] ), .YC(
        \CARRYB[10][5] ), .YS(\SUMB[10][5] ) );
  FAX1 S3_9_6 ( .A(n40), .B(\CARRYB[8][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[9][6] ), .YS(\SUMB[9][6] ) );
  FAX1 S2_9_5 ( .A(n39), .B(\CARRYB[8][5] ), .C(\SUMB[8][6] ), .YC(
        \CARRYB[9][5] ), .YS(\SUMB[9][5] ) );
  FAX1 S3_8_6 ( .A(n40), .B(\CARRYB[7][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[8][6] ), .YS(\SUMB[8][6] ) );
  FAX1 S2_8_5 ( .A(n39), .B(\CARRYB[7][5] ), .C(\SUMB[7][6] ), .YC(
        \CARRYB[8][5] ), .YS(\SUMB[8][5] ) );
  FAX1 S3_7_6 ( .A(n40), .B(\CARRYB[6][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S2_7_5 ( .A(n39), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S3_6_6 ( .A(n40), .B(\CARRYB[5][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_5 ( .A(n39), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S3_5_6 ( .A(n40), .B(\CARRYB[4][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_5 ( .A(n39), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S3_4_6 ( .A(n40), .B(\CARRYB[3][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_5 ( .A(n39), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S3_3_6 ( .A(n40), .B(\CARRYB[2][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  AND2X2 U9 ( .A(B[7]), .B(A[9]), .Y(\ab[9][7] ) );
  FAX1 S2_3_5 ( .A(n39), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S3_2_6 ( .A(n40), .B(n4), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), .YS(
        \SUMB[2][6] ) );
  NAND2X1 U10 ( .A(B[6]), .B(A[9]), .Y(n10) );
  FAX1 S2_2_5 ( .A(n39), .B(n3), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), .YS(
        \SUMB[2][5] ) );
  NAND2X1 U12 ( .A(B[5]), .B(A[9]), .Y(n12) );
  INVX4 U11 ( .A(n10), .Y(n40) );
  INVX4 U13 ( .A(n12), .Y(n39) );
  INVX4 U15 ( .A(n14), .Y(n38) );
  INVX4 U17 ( .A(n16), .Y(n37) );
  INVX4 U19 ( .A(n18), .Y(n36) );
  INVX4 U21 ( .A(n20), .Y(n35) );
  INVX4 U23 ( .A(n22), .Y(n34) );
  INVX2 U31 ( .A(A[0]), .Y(n41) );
  INVX2 U32 ( .A(A[1]), .Y(n42) );
  INVX2 U33 ( .A(B[0]), .Y(n43) );
  INVX2 U34 ( .A(B[1]), .Y(n44) );
  INVX2 U35 ( .A(B[2]), .Y(n45) );
  INVX2 U36 ( .A(B[3]), .Y(n46) );
  INVX2 U37 ( .A(B[4]), .Y(n47) );
  INVX2 U38 ( .A(B[5]), .Y(n48) );
  INVX2 U39 ( .A(B[6]), .Y(n49) );
  INVX2 U40 ( .A(B[7]), .Y(n50) );
endmodule


module CannyEdge_DW02_mult_14 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n35), .B(\SUMB[6][4] ), .Y(n3) );
  AND2X2 U3 ( .A(n32), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n36), .B(\SUMB[2][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n37), .B(\SUMB[2][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[2][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n39), .B(\SUMB[2][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n40), .B(\SUMB[2][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n41), .B(\SUMB[2][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n27), .B(\SUMB[4][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n33), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n11), .B(n43), .Y(n14) );
  AND2X2 U14 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n4), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[3][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][5] ), .Y(n27) );
  AND2X2 U27 ( .A(n23), .B(\SUMB[4][1] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][2] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][3] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][4] ), .Y(n31) );
  AND2X2 U31 ( .A(n28), .B(\SUMB[5][1] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][2] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][3] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][4] ), .Y(n35) );
  AND2X2 U35 ( .A(n21), .B(\SUMB[1][1] ), .Y(n36) );
  AND2X2 U36 ( .A(n15), .B(\SUMB[1][2] ), .Y(n37) );
  AND2X2 U37 ( .A(n16), .B(\SUMB[1][3] ), .Y(n38) );
  AND2X2 U38 ( .A(n17), .B(\SUMB[1][4] ), .Y(n39) );
  AND2X2 U39 ( .A(n18), .B(\SUMB[1][5] ), .Y(n40) );
  AND2X2 U40 ( .A(n19), .B(\SUMB[1][6] ), .Y(n41) );
  AND2X2 U41 ( .A(n20), .B(\ab[1][7] ), .Y(n42) );
  AND2X2 U42 ( .A(n10), .B(n42), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n13), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n12), .Y(n45) );
  XNOR2X1 U45 ( .A(n61), .B(n22), .Y(PRODUCT[9]) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n14), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n14), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n21), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n15), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n16), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n17), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n18), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n19), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n20), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n36), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n37), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n38), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n39), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n40), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n41), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n5), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n6), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n7), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n8), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n9), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n42), .B(n10), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n23), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n24), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n25), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n26), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n27), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n28), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n29), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n30), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n31), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n43), .B(n11), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n32), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n33), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n34), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n35), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n45), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n45), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n44), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n44), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n22), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_15 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [7:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , n9, n8, n7, n6, n5, n4, n3, n24, n22, n20,
         n18, n16, n14, n12, n10, \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[30][1] ,
         \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] ,
         \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[30][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] ,
         \CARRYB[28][1] , \CARRYB[28][0] , \CARRYB[27][3] , \CARRYB[27][2] ,
         \CARRYB[27][1] , \CARRYB[27][0] , \CARRYB[26][4] , \CARRYB[26][3] ,
         \CARRYB[26][2] , \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] ,
         \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][6] ,
         \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] ,
         \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][6] ,
         \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] ,
         \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] ,
         \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][6] ,
         \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] ,
         \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , n26, n27, n28, n29, n30, n31, n32,
         n33;

  XOR2X1 U31 ( .A(n33), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  AND2X1 U32 ( .A(B[7]), .B(A[0]), .Y(\ab[0][7] ) );
  AND2X1 U33 ( .A(B[6]), .B(A[0]), .Y(\ab[0][6] ) );
  AND2X1 U34 ( .A(B[5]), .B(A[0]), .Y(\ab[0][5] ) );
  AND2X1 U35 ( .A(B[4]), .B(A[0]), .Y(\ab[0][4] ) );
  AND2X1 U36 ( .A(B[3]), .B(A[0]), .Y(\ab[0][3] ) );
  AND2X1 U37 ( .A(B[2]), .B(A[0]), .Y(\ab[0][2] ) );
  AND2X1 U38 ( .A(B[1]), .B(A[0]), .Y(\ab[0][1] ) );
  AND2X1 U39 ( .A(B[0]), .B(A[0]), .Y(PRODUCT[0]) );
  FAX1 S4_0 ( .A(n33), .B(\CARRYB[30][0] ), .C(\SUMB[30][1] ), .YS(PRODUCT[31]) );
  FAX1 S1_30_0 ( .A(n33), .B(\CARRYB[29][0] ), .C(\SUMB[29][1] ), .YC(
        \CARRYB[30][0] ), .YS(PRODUCT[30]) );
  FAX1 S1_29_0 ( .A(n33), .B(\CARRYB[28][0] ), .C(\SUMB[28][1] ), .YC(
        \CARRYB[29][0] ), .YS(PRODUCT[29]) );
  FAX1 S1_28_0 ( .A(n33), .B(\CARRYB[27][0] ), .C(\SUMB[27][1] ), .YC(
        \CARRYB[28][0] ), .YS(PRODUCT[28]) );
  FAX1 S1_27_0 ( .A(n33), .B(\CARRYB[26][0] ), .C(\SUMB[26][1] ), .YC(
        \CARRYB[27][0] ), .YS(PRODUCT[27]) );
  FAX1 S1_26_0 ( .A(n33), .B(\CARRYB[25][0] ), .C(\SUMB[25][1] ), .YC(
        \CARRYB[26][0] ), .YS(PRODUCT[26]) );
  FAX1 S1_25_0 ( .A(n33), .B(\CARRYB[24][0] ), .C(\SUMB[24][1] ), .YC(
        \CARRYB[25][0] ), .YS(PRODUCT[25]) );
  FAX1 S1_24_0 ( .A(n33), .B(\CARRYB[23][0] ), .C(\SUMB[23][1] ), .YC(
        \CARRYB[24][0] ), .YS(PRODUCT[24]) );
  FAX1 S1_23_0 ( .A(n33), .B(\CARRYB[22][0] ), .C(\SUMB[22][1] ), .YC(
        \CARRYB[23][0] ), .YS(PRODUCT[23]) );
  FAX1 S1_22_0 ( .A(n33), .B(\CARRYB[21][0] ), .C(\SUMB[21][1] ), .YC(
        \CARRYB[22][0] ), .YS(PRODUCT[22]) );
  FAX1 S1_21_0 ( .A(n33), .B(\CARRYB[20][0] ), .C(\SUMB[20][1] ), .YC(
        \CARRYB[21][0] ), .YS(PRODUCT[21]) );
  FAX1 S1_20_0 ( .A(n33), .B(\CARRYB[19][0] ), .C(\SUMB[19][1] ), .YC(
        \CARRYB[20][0] ), .YS(PRODUCT[20]) );
  FAX1 S1_19_0 ( .A(n33), .B(\CARRYB[18][0] ), .C(\SUMB[18][1] ), .YC(
        \CARRYB[19][0] ), .YS(PRODUCT[19]) );
  FAX1 S1_18_0 ( .A(n33), .B(\CARRYB[17][0] ), .C(\SUMB[17][1] ), .YC(
        \CARRYB[18][0] ), .YS(PRODUCT[18]) );
  FAX1 S1_17_0 ( .A(n33), .B(\CARRYB[16][0] ), .C(\SUMB[16][1] ), .YC(
        \CARRYB[17][0] ), .YS(PRODUCT[17]) );
  FAX1 S1_16_0 ( .A(n33), .B(\CARRYB[15][0] ), .C(\SUMB[15][1] ), .YC(
        \CARRYB[16][0] ), .YS(PRODUCT[16]) );
  FAX1 S1_15_0 ( .A(n33), .B(\CARRYB[14][0] ), .C(\SUMB[14][1] ), .YC(
        \CARRYB[15][0] ), .YS(PRODUCT[15]) );
  FAX1 S1_14_0 ( .A(n33), .B(\CARRYB[13][0] ), .C(\SUMB[13][1] ), .YC(
        \CARRYB[14][0] ), .YS(PRODUCT[14]) );
  FAX1 S1_13_0 ( .A(n33), .B(\CARRYB[12][0] ), .C(\SUMB[12][1] ), .YC(
        \CARRYB[13][0] ), .YS(PRODUCT[13]) );
  FAX1 S1_12_0 ( .A(n33), .B(\CARRYB[11][0] ), .C(\SUMB[11][1] ), .YC(
        \CARRYB[12][0] ), .YS(PRODUCT[12]) );
  FAX1 S1_11_0 ( .A(n33), .B(\CARRYB[10][0] ), .C(\SUMB[10][1] ), .YC(
        \CARRYB[11][0] ), .YS(PRODUCT[11]) );
  FAX1 S1_10_0 ( .A(n33), .B(\CARRYB[9][0] ), .C(\SUMB[9][1] ), .YC(
        \CARRYB[10][0] ), .YS(PRODUCT[10]) );
  FAX1 S1_9_0 ( .A(n33), .B(\CARRYB[8][0] ), .C(\SUMB[8][1] ), .YC(
        \CARRYB[9][0] ), .YS(PRODUCT[9]) );
  FAX1 S1_8_0 ( .A(n33), .B(\CARRYB[7][0] ), .C(\SUMB[7][1] ), .YC(
        \CARRYB[8][0] ), .YS(PRODUCT[8]) );
  FAX1 S1_7_0 ( .A(n33), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(PRODUCT[7]) );
  FAX1 S1_6_0 ( .A(n33), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(PRODUCT[6]) );
  FAX1 S1_5_0 ( .A(n33), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(PRODUCT[5]) );
  FAX1 S1_4_0 ( .A(n33), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(PRODUCT[4]) );
  FAX1 S1_3_0 ( .A(n33), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(PRODUCT[3]) );
  FAX1 S1_2_0 ( .A(n33), .B(n3), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), .YS(
        PRODUCT[2]) );
  XOR2X1 U30 ( .A(n26), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  AND2X2 U2 ( .A(\ab[0][1] ), .B(n33), .Y(n3) );
  NAND2X1 U23 ( .A(B[0]), .B(A[9]), .Y(n24) );
  FAX1 S2_30_1 ( .A(n26), .B(\CARRYB[29][1] ), .C(\SUMB[29][2] ), .YS(
        \SUMB[30][1] ) );
  FAX1 S2_29_1 ( .A(n26), .B(\CARRYB[28][1] ), .C(\SUMB[28][2] ), .YC(
        \CARRYB[29][1] ), .YS(\SUMB[29][1] ) );
  FAX1 S2_28_1 ( .A(n26), .B(\CARRYB[27][1] ), .C(\SUMB[27][2] ), .YC(
        \CARRYB[28][1] ), .YS(\SUMB[28][1] ) );
  FAX1 S2_27_1 ( .A(n26), .B(\CARRYB[26][1] ), .C(\SUMB[26][2] ), .YC(
        \CARRYB[27][1] ), .YS(\SUMB[27][1] ) );
  FAX1 S2_26_1 ( .A(n26), .B(\CARRYB[25][1] ), .C(\SUMB[25][2] ), .YC(
        \CARRYB[26][1] ), .YS(\SUMB[26][1] ) );
  FAX1 S2_25_1 ( .A(n26), .B(\CARRYB[24][1] ), .C(\SUMB[24][2] ), .YC(
        \CARRYB[25][1] ), .YS(\SUMB[25][1] ) );
  FAX1 S2_24_1 ( .A(n26), .B(\CARRYB[23][1] ), .C(\SUMB[23][2] ), .YC(
        \CARRYB[24][1] ), .YS(\SUMB[24][1] ) );
  FAX1 S2_23_1 ( .A(n26), .B(\CARRYB[22][1] ), .C(\SUMB[22][2] ), .YC(
        \CARRYB[23][1] ), .YS(\SUMB[23][1] ) );
  FAX1 S2_22_1 ( .A(n26), .B(\CARRYB[21][1] ), .C(\SUMB[21][2] ), .YC(
        \CARRYB[22][1] ), .YS(\SUMB[22][1] ) );
  FAX1 S2_21_1 ( .A(n26), .B(\CARRYB[20][1] ), .C(\SUMB[20][2] ), .YC(
        \CARRYB[21][1] ), .YS(\SUMB[21][1] ) );
  FAX1 S2_20_1 ( .A(n26), .B(\CARRYB[19][1] ), .C(\SUMB[19][2] ), .YC(
        \CARRYB[20][1] ), .YS(\SUMB[20][1] ) );
  FAX1 S2_19_1 ( .A(n26), .B(\CARRYB[18][1] ), .C(\SUMB[18][2] ), .YC(
        \CARRYB[19][1] ), .YS(\SUMB[19][1] ) );
  FAX1 S2_18_1 ( .A(n26), .B(\CARRYB[17][1] ), .C(\SUMB[17][2] ), .YC(
        \CARRYB[18][1] ), .YS(\SUMB[18][1] ) );
  FAX1 S2_17_1 ( .A(n26), .B(\CARRYB[16][1] ), .C(\SUMB[16][2] ), .YC(
        \CARRYB[17][1] ), .YS(\SUMB[17][1] ) );
  FAX1 S2_16_1 ( .A(n26), .B(\CARRYB[15][1] ), .C(\SUMB[15][2] ), .YC(
        \CARRYB[16][1] ), .YS(\SUMB[16][1] ) );
  FAX1 S2_15_1 ( .A(n26), .B(\CARRYB[14][1] ), .C(\SUMB[14][2] ), .YC(
        \CARRYB[15][1] ), .YS(\SUMB[15][1] ) );
  FAX1 S2_14_1 ( .A(n26), .B(\CARRYB[13][1] ), .C(\SUMB[13][2] ), .YC(
        \CARRYB[14][1] ), .YS(\SUMB[14][1] ) );
  FAX1 S2_13_1 ( .A(n26), .B(\CARRYB[12][1] ), .C(\SUMB[12][2] ), .YC(
        \CARRYB[13][1] ), .YS(\SUMB[13][1] ) );
  FAX1 S2_12_1 ( .A(n26), .B(\CARRYB[11][1] ), .C(\SUMB[11][2] ), .YC(
        \CARRYB[12][1] ), .YS(\SUMB[12][1] ) );
  FAX1 S2_11_1 ( .A(n26), .B(\CARRYB[10][1] ), .C(\SUMB[10][2] ), .YC(
        \CARRYB[11][1] ), .YS(\SUMB[11][1] ) );
  FAX1 S2_10_1 ( .A(n26), .B(\CARRYB[9][1] ), .C(\SUMB[9][2] ), .YC(
        \CARRYB[10][1] ), .YS(\SUMB[10][1] ) );
  FAX1 S2_9_1 ( .A(n26), .B(\CARRYB[8][1] ), .C(\SUMB[8][2] ), .YC(
        \CARRYB[9][1] ), .YS(\SUMB[9][1] ) );
  FAX1 S2_8_1 ( .A(n26), .B(\CARRYB[7][1] ), .C(\SUMB[7][2] ), .YC(
        \CARRYB[8][1] ), .YS(\SUMB[8][1] ) );
  FAX1 S2_7_1 ( .A(n26), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S2_6_1 ( .A(n26), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_5_1 ( .A(n26), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_4_1 ( .A(n26), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_3_1 ( .A(n26), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_2_1 ( .A(n26), .B(n4), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), .YS(
        \SUMB[2][1] ) );
  XOR2X1 U29 ( .A(n27), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  AND2X2 U3 ( .A(\ab[0][2] ), .B(n26), .Y(n4) );
  NAND2X1 U21 ( .A(B[1]), .B(A[9]), .Y(n22) );
  FAX1 S2_29_2 ( .A(n27), .B(\CARRYB[28][2] ), .C(\SUMB[28][3] ), .YS(
        \SUMB[29][2] ) );
  FAX1 S2_28_2 ( .A(n27), .B(\CARRYB[27][2] ), .C(\SUMB[27][3] ), .YC(
        \CARRYB[28][2] ), .YS(\SUMB[28][2] ) );
  FAX1 S2_27_2 ( .A(n27), .B(\CARRYB[26][2] ), .C(\SUMB[26][3] ), .YC(
        \CARRYB[27][2] ), .YS(\SUMB[27][2] ) );
  FAX1 S2_26_2 ( .A(n27), .B(\CARRYB[25][2] ), .C(\SUMB[25][3] ), .YC(
        \CARRYB[26][2] ), .YS(\SUMB[26][2] ) );
  FAX1 S2_25_2 ( .A(n27), .B(\CARRYB[24][2] ), .C(\SUMB[24][3] ), .YC(
        \CARRYB[25][2] ), .YS(\SUMB[25][2] ) );
  FAX1 S2_24_2 ( .A(n27), .B(\CARRYB[23][2] ), .C(\SUMB[23][3] ), .YC(
        \CARRYB[24][2] ), .YS(\SUMB[24][2] ) );
  FAX1 S2_23_2 ( .A(n27), .B(\CARRYB[22][2] ), .C(\SUMB[22][3] ), .YC(
        \CARRYB[23][2] ), .YS(\SUMB[23][2] ) );
  FAX1 S2_22_2 ( .A(n27), .B(\CARRYB[21][2] ), .C(\SUMB[21][3] ), .YC(
        \CARRYB[22][2] ), .YS(\SUMB[22][2] ) );
  FAX1 S2_21_2 ( .A(n27), .B(\CARRYB[20][2] ), .C(\SUMB[20][3] ), .YC(
        \CARRYB[21][2] ), .YS(\SUMB[21][2] ) );
  FAX1 S2_20_2 ( .A(n27), .B(\CARRYB[19][2] ), .C(\SUMB[19][3] ), .YC(
        \CARRYB[20][2] ), .YS(\SUMB[20][2] ) );
  FAX1 S2_19_2 ( .A(n27), .B(\CARRYB[18][2] ), .C(\SUMB[18][3] ), .YC(
        \CARRYB[19][2] ), .YS(\SUMB[19][2] ) );
  FAX1 S2_18_2 ( .A(n27), .B(\CARRYB[17][2] ), .C(\SUMB[17][3] ), .YC(
        \CARRYB[18][2] ), .YS(\SUMB[18][2] ) );
  FAX1 S2_17_2 ( .A(n27), .B(\CARRYB[16][2] ), .C(\SUMB[16][3] ), .YC(
        \CARRYB[17][2] ), .YS(\SUMB[17][2] ) );
  FAX1 S2_16_2 ( .A(n27), .B(\CARRYB[15][2] ), .C(\SUMB[15][3] ), .YC(
        \CARRYB[16][2] ), .YS(\SUMB[16][2] ) );
  FAX1 S2_15_2 ( .A(n27), .B(\CARRYB[14][2] ), .C(\SUMB[14][3] ), .YC(
        \CARRYB[15][2] ), .YS(\SUMB[15][2] ) );
  FAX1 S2_14_2 ( .A(n27), .B(\CARRYB[13][2] ), .C(\SUMB[13][3] ), .YC(
        \CARRYB[14][2] ), .YS(\SUMB[14][2] ) );
  FAX1 S2_13_2 ( .A(n27), .B(\CARRYB[12][2] ), .C(\SUMB[12][3] ), .YC(
        \CARRYB[13][2] ), .YS(\SUMB[13][2] ) );
  FAX1 S2_12_2 ( .A(n27), .B(\CARRYB[11][2] ), .C(\SUMB[11][3] ), .YC(
        \CARRYB[12][2] ), .YS(\SUMB[12][2] ) );
  FAX1 S2_11_2 ( .A(n27), .B(\CARRYB[10][2] ), .C(\SUMB[10][3] ), .YC(
        \CARRYB[11][2] ), .YS(\SUMB[11][2] ) );
  FAX1 S2_10_2 ( .A(n27), .B(\CARRYB[9][2] ), .C(\SUMB[9][3] ), .YC(
        \CARRYB[10][2] ), .YS(\SUMB[10][2] ) );
  FAX1 S2_9_2 ( .A(n27), .B(\CARRYB[8][2] ), .C(\SUMB[8][3] ), .YC(
        \CARRYB[9][2] ), .YS(\SUMB[9][2] ) );
  FAX1 S2_8_2 ( .A(n27), .B(\CARRYB[7][2] ), .C(\SUMB[7][3] ), .YC(
        \CARRYB[8][2] ), .YS(\SUMB[8][2] ) );
  FAX1 S2_7_2 ( .A(n27), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(n27), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_5_2 ( .A(n27), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_4_2 ( .A(n27), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_3_2 ( .A(n27), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_2_2 ( .A(n27), .B(n5), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), .YS(
        \SUMB[2][2] ) );
  XOR2X1 U28 ( .A(n29), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  AND2X2 U4 ( .A(\ab[0][3] ), .B(n27), .Y(n5) );
  NAND2X1 U19 ( .A(B[2]), .B(A[9]), .Y(n20) );
  FAX1 S2_28_3 ( .A(n29), .B(\CARRYB[27][3] ), .C(\SUMB[27][4] ), .YS(
        \SUMB[28][3] ) );
  FAX1 S2_27_3 ( .A(n29), .B(\CARRYB[26][3] ), .C(\SUMB[26][4] ), .YC(
        \CARRYB[27][3] ), .YS(\SUMB[27][3] ) );
  FAX1 S2_26_3 ( .A(n29), .B(\CARRYB[25][3] ), .C(\SUMB[25][4] ), .YC(
        \CARRYB[26][3] ), .YS(\SUMB[26][3] ) );
  FAX1 S2_25_3 ( .A(n29), .B(\CARRYB[24][3] ), .C(\SUMB[24][4] ), .YC(
        \CARRYB[25][3] ), .YS(\SUMB[25][3] ) );
  FAX1 S2_24_3 ( .A(n29), .B(\CARRYB[23][3] ), .C(\SUMB[23][4] ), .YC(
        \CARRYB[24][3] ), .YS(\SUMB[24][3] ) );
  FAX1 S2_23_3 ( .A(n29), .B(\CARRYB[22][3] ), .C(\SUMB[22][4] ), .YC(
        \CARRYB[23][3] ), .YS(\SUMB[23][3] ) );
  FAX1 S2_22_3 ( .A(n29), .B(\CARRYB[21][3] ), .C(\SUMB[21][4] ), .YC(
        \CARRYB[22][3] ), .YS(\SUMB[22][3] ) );
  FAX1 S2_21_3 ( .A(n29), .B(\CARRYB[20][3] ), .C(\SUMB[20][4] ), .YC(
        \CARRYB[21][3] ), .YS(\SUMB[21][3] ) );
  FAX1 S2_20_3 ( .A(n29), .B(\CARRYB[19][3] ), .C(\SUMB[19][4] ), .YC(
        \CARRYB[20][3] ), .YS(\SUMB[20][3] ) );
  FAX1 S2_19_3 ( .A(n29), .B(\CARRYB[18][3] ), .C(\SUMB[18][4] ), .YC(
        \CARRYB[19][3] ), .YS(\SUMB[19][3] ) );
  FAX1 S2_18_3 ( .A(n29), .B(\CARRYB[17][3] ), .C(\SUMB[17][4] ), .YC(
        \CARRYB[18][3] ), .YS(\SUMB[18][3] ) );
  FAX1 S2_17_3 ( .A(n29), .B(\CARRYB[16][3] ), .C(\SUMB[16][4] ), .YC(
        \CARRYB[17][3] ), .YS(\SUMB[17][3] ) );
  FAX1 S2_16_3 ( .A(n29), .B(\CARRYB[15][3] ), .C(\SUMB[15][4] ), .YC(
        \CARRYB[16][3] ), .YS(\SUMB[16][3] ) );
  FAX1 S2_15_3 ( .A(n29), .B(\CARRYB[14][3] ), .C(\SUMB[14][4] ), .YC(
        \CARRYB[15][3] ), .YS(\SUMB[15][3] ) );
  FAX1 S2_14_3 ( .A(n29), .B(\CARRYB[13][3] ), .C(\SUMB[13][4] ), .YC(
        \CARRYB[14][3] ), .YS(\SUMB[14][3] ) );
  FAX1 S2_13_3 ( .A(n29), .B(\CARRYB[12][3] ), .C(\SUMB[12][4] ), .YC(
        \CARRYB[13][3] ), .YS(\SUMB[13][3] ) );
  FAX1 S2_12_3 ( .A(n29), .B(\CARRYB[11][3] ), .C(\SUMB[11][4] ), .YC(
        \CARRYB[12][3] ), .YS(\SUMB[12][3] ) );
  FAX1 S2_11_3 ( .A(n29), .B(\CARRYB[10][3] ), .C(\SUMB[10][4] ), .YC(
        \CARRYB[11][3] ), .YS(\SUMB[11][3] ) );
  FAX1 S2_10_3 ( .A(n29), .B(\CARRYB[9][3] ), .C(\SUMB[9][4] ), .YC(
        \CARRYB[10][3] ), .YS(\SUMB[10][3] ) );
  FAX1 S2_9_3 ( .A(n29), .B(\CARRYB[8][3] ), .C(\SUMB[8][4] ), .YC(
        \CARRYB[9][3] ), .YS(\SUMB[9][3] ) );
  FAX1 S2_8_3 ( .A(n29), .B(\CARRYB[7][3] ), .C(\SUMB[7][4] ), .YC(
        \CARRYB[8][3] ), .YS(\SUMB[8][3] ) );
  FAX1 S2_7_3 ( .A(n29), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(n29), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(n29), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_4_3 ( .A(n29), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_3_3 ( .A(n29), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_2_3 ( .A(n29), .B(n6), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), .YS(
        \SUMB[2][3] ) );
  XOR2X1 U27 ( .A(n28), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  AND2X2 U5 ( .A(\ab[0][4] ), .B(n29), .Y(n6) );
  NAND2X1 U15 ( .A(B[3]), .B(A[9]), .Y(n16) );
  FAX1 S2_27_4 ( .A(n28), .B(\CARRYB[26][4] ), .C(\SUMB[26][5] ), .YS(
        \SUMB[27][4] ) );
  FAX1 S2_26_4 ( .A(n28), .B(\CARRYB[25][4] ), .C(\SUMB[25][5] ), .YC(
        \CARRYB[26][4] ), .YS(\SUMB[26][4] ) );
  FAX1 S2_25_4 ( .A(n28), .B(\CARRYB[24][4] ), .C(\SUMB[24][5] ), .YC(
        \CARRYB[25][4] ), .YS(\SUMB[25][4] ) );
  FAX1 S2_24_4 ( .A(n28), .B(\CARRYB[23][4] ), .C(\SUMB[23][5] ), .YC(
        \CARRYB[24][4] ), .YS(\SUMB[24][4] ) );
  FAX1 S2_23_4 ( .A(n28), .B(\CARRYB[22][4] ), .C(\SUMB[22][5] ), .YC(
        \CARRYB[23][4] ), .YS(\SUMB[23][4] ) );
  FAX1 S2_22_4 ( .A(n28), .B(\CARRYB[21][4] ), .C(\SUMB[21][5] ), .YC(
        \CARRYB[22][4] ), .YS(\SUMB[22][4] ) );
  FAX1 S2_21_4 ( .A(n28), .B(\CARRYB[20][4] ), .C(\SUMB[20][5] ), .YC(
        \CARRYB[21][4] ), .YS(\SUMB[21][4] ) );
  FAX1 S2_20_4 ( .A(n28), .B(\CARRYB[19][4] ), .C(\SUMB[19][5] ), .YC(
        \CARRYB[20][4] ), .YS(\SUMB[20][4] ) );
  FAX1 S2_19_4 ( .A(n28), .B(\CARRYB[18][4] ), .C(\SUMB[18][5] ), .YC(
        \CARRYB[19][4] ), .YS(\SUMB[19][4] ) );
  FAX1 S2_18_4 ( .A(n28), .B(\CARRYB[17][4] ), .C(\SUMB[17][5] ), .YC(
        \CARRYB[18][4] ), .YS(\SUMB[18][4] ) );
  FAX1 S2_17_4 ( .A(n28), .B(\CARRYB[16][4] ), .C(\SUMB[16][5] ), .YC(
        \CARRYB[17][4] ), .YS(\SUMB[17][4] ) );
  FAX1 S2_16_4 ( .A(n28), .B(\CARRYB[15][4] ), .C(\SUMB[15][5] ), .YC(
        \CARRYB[16][4] ), .YS(\SUMB[16][4] ) );
  FAX1 S2_15_4 ( .A(n28), .B(\CARRYB[14][4] ), .C(\SUMB[14][5] ), .YC(
        \CARRYB[15][4] ), .YS(\SUMB[15][4] ) );
  FAX1 S2_14_4 ( .A(n28), .B(\CARRYB[13][4] ), .C(\SUMB[13][5] ), .YC(
        \CARRYB[14][4] ), .YS(\SUMB[14][4] ) );
  FAX1 S2_13_4 ( .A(n28), .B(\CARRYB[12][4] ), .C(\SUMB[12][5] ), .YC(
        \CARRYB[13][4] ), .YS(\SUMB[13][4] ) );
  FAX1 S2_12_4 ( .A(n28), .B(\CARRYB[11][4] ), .C(\SUMB[11][5] ), .YC(
        \CARRYB[12][4] ), .YS(\SUMB[12][4] ) );
  FAX1 S2_11_4 ( .A(n28), .B(\CARRYB[10][4] ), .C(\SUMB[10][5] ), .YC(
        \CARRYB[11][4] ), .YS(\SUMB[11][4] ) );
  FAX1 S2_10_4 ( .A(n28), .B(\CARRYB[9][4] ), .C(\SUMB[9][5] ), .YC(
        \CARRYB[10][4] ), .YS(\SUMB[10][4] ) );
  FAX1 S2_9_4 ( .A(n28), .B(\CARRYB[8][4] ), .C(\SUMB[8][5] ), .YC(
        \CARRYB[9][4] ), .YS(\SUMB[9][4] ) );
  FAX1 S2_8_4 ( .A(n28), .B(\CARRYB[7][4] ), .C(\SUMB[7][5] ), .YC(
        \CARRYB[8][4] ), .YS(\SUMB[8][4] ) );
  FAX1 S2_7_4 ( .A(n28), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(n28), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(n28), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(n28), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_3_4 ( .A(n28), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_2_4 ( .A(n28), .B(n7), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), .YS(
        \SUMB[2][4] ) );
  XOR2X1 U26 ( .A(n30), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  AND2X2 U6 ( .A(\ab[0][5] ), .B(n28), .Y(n7) );
  NAND2X1 U17 ( .A(B[4]), .B(A[9]), .Y(n18) );
  FAX1 S2_26_5 ( .A(n30), .B(\CARRYB[25][5] ), .C(\SUMB[25][6] ), .YS(
        \SUMB[26][5] ) );
  FAX1 S3_25_6 ( .A(n31), .B(\CARRYB[24][6] ), .C(n32), .YS(\SUMB[25][6] ) );
  FAX1 S2_25_5 ( .A(n30), .B(\CARRYB[24][5] ), .C(\SUMB[24][6] ), .YC(
        \CARRYB[25][5] ), .YS(\SUMB[25][5] ) );
  FAX1 S3_24_6 ( .A(n31), .B(\CARRYB[23][6] ), .C(n32), .YC(\CARRYB[24][6] ), 
        .YS(\SUMB[24][6] ) );
  FAX1 S2_24_5 ( .A(n30), .B(\CARRYB[23][5] ), .C(\SUMB[23][6] ), .YC(
        \CARRYB[24][5] ), .YS(\SUMB[24][5] ) );
  FAX1 S3_23_6 ( .A(n31), .B(\CARRYB[22][6] ), .C(n32), .YC(\CARRYB[23][6] ), 
        .YS(\SUMB[23][6] ) );
  FAX1 S2_23_5 ( .A(n30), .B(\CARRYB[22][5] ), .C(\SUMB[22][6] ), .YC(
        \CARRYB[23][5] ), .YS(\SUMB[23][5] ) );
  FAX1 S3_22_6 ( .A(n31), .B(\CARRYB[21][6] ), .C(n32), .YC(\CARRYB[22][6] ), 
        .YS(\SUMB[22][6] ) );
  FAX1 S2_22_5 ( .A(n30), .B(\CARRYB[21][5] ), .C(\SUMB[21][6] ), .YC(
        \CARRYB[22][5] ), .YS(\SUMB[22][5] ) );
  FAX1 S3_21_6 ( .A(n31), .B(\CARRYB[20][6] ), .C(n32), .YC(\CARRYB[21][6] ), 
        .YS(\SUMB[21][6] ) );
  FAX1 S2_21_5 ( .A(n30), .B(\CARRYB[20][5] ), .C(\SUMB[20][6] ), .YC(
        \CARRYB[21][5] ), .YS(\SUMB[21][5] ) );
  FAX1 S3_20_6 ( .A(n31), .B(\CARRYB[19][6] ), .C(n32), .YC(\CARRYB[20][6] ), 
        .YS(\SUMB[20][6] ) );
  FAX1 S2_20_5 ( .A(n30), .B(\CARRYB[19][5] ), .C(\SUMB[19][6] ), .YC(
        \CARRYB[20][5] ), .YS(\SUMB[20][5] ) );
  FAX1 S3_19_6 ( .A(n31), .B(\CARRYB[18][6] ), .C(n32), .YC(\CARRYB[19][6] ), 
        .YS(\SUMB[19][6] ) );
  FAX1 S2_19_5 ( .A(n30), .B(\CARRYB[18][5] ), .C(\SUMB[18][6] ), .YC(
        \CARRYB[19][5] ), .YS(\SUMB[19][5] ) );
  FAX1 S3_18_6 ( .A(n31), .B(\CARRYB[17][6] ), .C(n32), .YC(\CARRYB[18][6] ), 
        .YS(\SUMB[18][6] ) );
  FAX1 S2_18_5 ( .A(n30), .B(\CARRYB[17][5] ), .C(\SUMB[17][6] ), .YC(
        \CARRYB[18][5] ), .YS(\SUMB[18][5] ) );
  FAX1 S3_17_6 ( .A(n31), .B(\CARRYB[16][6] ), .C(n32), .YC(\CARRYB[17][6] ), 
        .YS(\SUMB[17][6] ) );
  FAX1 S2_17_5 ( .A(n30), .B(\CARRYB[16][5] ), .C(\SUMB[16][6] ), .YC(
        \CARRYB[17][5] ), .YS(\SUMB[17][5] ) );
  FAX1 S3_16_6 ( .A(n31), .B(\CARRYB[15][6] ), .C(n32), .YC(\CARRYB[16][6] ), 
        .YS(\SUMB[16][6] ) );
  FAX1 S2_16_5 ( .A(n30), .B(\CARRYB[15][5] ), .C(\SUMB[15][6] ), .YC(
        \CARRYB[16][5] ), .YS(\SUMB[16][5] ) );
  FAX1 S3_15_6 ( .A(n31), .B(\CARRYB[14][6] ), .C(n32), .YC(\CARRYB[15][6] ), 
        .YS(\SUMB[15][6] ) );
  FAX1 S2_15_5 ( .A(n30), .B(\CARRYB[14][5] ), .C(\SUMB[14][6] ), .YC(
        \CARRYB[15][5] ), .YS(\SUMB[15][5] ) );
  FAX1 S3_14_6 ( .A(n31), .B(\CARRYB[13][6] ), .C(n32), .YC(\CARRYB[14][6] ), 
        .YS(\SUMB[14][6] ) );
  FAX1 S2_14_5 ( .A(n30), .B(\CARRYB[13][5] ), .C(\SUMB[13][6] ), .YC(
        \CARRYB[14][5] ), .YS(\SUMB[14][5] ) );
  FAX1 S3_13_6 ( .A(n31), .B(\CARRYB[12][6] ), .C(n32), .YC(\CARRYB[13][6] ), 
        .YS(\SUMB[13][6] ) );
  FAX1 S2_13_5 ( .A(n30), .B(\CARRYB[12][5] ), .C(\SUMB[12][6] ), .YC(
        \CARRYB[13][5] ), .YS(\SUMB[13][5] ) );
  FAX1 S3_12_6 ( .A(n31), .B(\CARRYB[11][6] ), .C(n32), .YC(\CARRYB[12][6] ), 
        .YS(\SUMB[12][6] ) );
  FAX1 S2_12_5 ( .A(n30), .B(\CARRYB[11][5] ), .C(\SUMB[11][6] ), .YC(
        \CARRYB[12][5] ), .YS(\SUMB[12][5] ) );
  FAX1 S3_11_6 ( .A(n31), .B(\CARRYB[10][6] ), .C(n32), .YC(\CARRYB[11][6] ), 
        .YS(\SUMB[11][6] ) );
  FAX1 S2_11_5 ( .A(n30), .B(\CARRYB[10][5] ), .C(\SUMB[10][6] ), .YC(
        \CARRYB[11][5] ), .YS(\SUMB[11][5] ) );
  FAX1 S3_10_6 ( .A(n31), .B(\CARRYB[9][6] ), .C(n32), .YC(\CARRYB[10][6] ), 
        .YS(\SUMB[10][6] ) );
  FAX1 S2_10_5 ( .A(n30), .B(\CARRYB[9][5] ), .C(\SUMB[9][6] ), .YC(
        \CARRYB[10][5] ), .YS(\SUMB[10][5] ) );
  FAX1 S3_9_6 ( .A(n31), .B(\CARRYB[8][6] ), .C(n32), .YC(\CARRYB[9][6] ), 
        .YS(\SUMB[9][6] ) );
  FAX1 S2_9_5 ( .A(n30), .B(\CARRYB[8][5] ), .C(\SUMB[8][6] ), .YC(
        \CARRYB[9][5] ), .YS(\SUMB[9][5] ) );
  FAX1 S3_8_6 ( .A(n31), .B(\CARRYB[7][6] ), .C(n32), .YC(\CARRYB[8][6] ), 
        .YS(\SUMB[8][6] ) );
  FAX1 S2_8_5 ( .A(n30), .B(\CARRYB[7][5] ), .C(\SUMB[7][6] ), .YC(
        \CARRYB[8][5] ), .YS(\SUMB[8][5] ) );
  FAX1 S3_7_6 ( .A(n31), .B(\CARRYB[6][6] ), .C(n32), .YC(\CARRYB[7][6] ), 
        .YS(\SUMB[7][6] ) );
  FAX1 S2_7_5 ( .A(n30), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S3_6_6 ( .A(n31), .B(\CARRYB[5][6] ), .C(n32), .YC(\CARRYB[6][6] ), 
        .YS(\SUMB[6][6] ) );
  FAX1 S2_6_5 ( .A(n30), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S3_5_6 ( .A(n31), .B(\CARRYB[4][6] ), .C(n32), .YC(\CARRYB[5][6] ), 
        .YS(\SUMB[5][6] ) );
  FAX1 S2_5_5 ( .A(n30), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S3_4_6 ( .A(n31), .B(\CARRYB[3][6] ), .C(n32), .YC(\CARRYB[4][6] ), 
        .YS(\SUMB[4][6] ) );
  FAX1 S2_4_5 ( .A(n30), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S3_3_6 ( .A(n31), .B(\CARRYB[2][6] ), .C(n32), .YC(\CARRYB[3][6] ), 
        .YS(\SUMB[3][6] ) );
  FAX1 S2_3_5 ( .A(n30), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S3_2_6 ( .A(n31), .B(n9), .C(n32), .YC(\CARRYB[2][6] ), .YS(
        \SUMB[2][6] ) );
  NAND2X1 U9 ( .A(B[7]), .B(A[9]), .Y(n10) );
  AND2X2 U8 ( .A(\ab[0][7] ), .B(n31), .Y(n9) );
  FAX1 S2_2_5 ( .A(n30), .B(n8), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), .YS(
        \SUMB[2][5] ) );
  XOR2X1 U25 ( .A(n31), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  NAND2X1 U11 ( .A(B[6]), .B(A[9]), .Y(n12) );
  AND2X2 U7 ( .A(\ab[0][6] ), .B(n30), .Y(n8) );
  NAND2X1 U13 ( .A(B[5]), .B(A[9]), .Y(n14) );
  INVX4 U10 ( .A(n10), .Y(n32) );
  INVX4 U12 ( .A(n12), .Y(n31) );
  INVX4 U14 ( .A(n14), .Y(n30) );
  INVX4 U16 ( .A(n16), .Y(n29) );
  INVX4 U18 ( .A(n18), .Y(n28) );
  INVX4 U20 ( .A(n20), .Y(n27) );
  INVX4 U22 ( .A(n22), .Y(n26) );
  INVX4 U24 ( .A(n24), .Y(n33) );
endmodule


module CannyEdge_DW02_mult_16 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n22), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n21), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n20), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n18), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n17), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n16), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n73), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n33), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n34), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n35), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n36), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n37), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n38), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n39), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n33), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n34), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n35), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n36), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n37), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n38), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n39), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n77), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n75), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n72), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  NOR2X1 U114 ( .A(n83), .B(n82), .Y(\ab[2][7] ) );
  NOR2X1 U115 ( .A(n83), .B(n81), .Y(\ab[2][6] ) );
  NOR2X1 U116 ( .A(n83), .B(n80), .Y(\ab[2][5] ) );
  NOR2X1 U117 ( .A(n83), .B(n79), .Y(\ab[2][4] ) );
  NOR2X1 U118 ( .A(n83), .B(n78), .Y(\ab[2][3] ) );
  NOR2X1 U119 ( .A(n83), .B(n76), .Y(\ab[2][2] ) );
  NOR2X1 U120 ( .A(n83), .B(n74), .Y(\ab[2][1] ) );
  NOR2X1 U121 ( .A(n83), .B(n71), .Y(\ab[2][0] ) );
  NOR2X1 U122 ( .A(n82), .B(n84), .Y(\ab[1][7] ) );
  NOR2X1 U123 ( .A(n81), .B(n84), .Y(\ab[1][6] ) );
  NOR2X1 U124 ( .A(n80), .B(n84), .Y(\ab[1][5] ) );
  NOR2X1 U125 ( .A(n79), .B(n84), .Y(\ab[1][4] ) );
  NOR2X1 U126 ( .A(n78), .B(n84), .Y(\ab[1][3] ) );
  NOR2X1 U127 ( .A(n76), .B(n84), .Y(\ab[1][2] ) );
  NOR2X1 U128 ( .A(n74), .B(n84), .Y(\ab[1][1] ) );
  NOR2X1 U129 ( .A(n71), .B(n84), .Y(\ab[1][0] ) );
  NOR2X1 U130 ( .A(n82), .B(n85), .Y(\ab[0][7] ) );
  NOR2X1 U131 ( .A(n81), .B(n85), .Y(\ab[0][6] ) );
  NOR2X1 U132 ( .A(n80), .B(n85), .Y(\ab[0][5] ) );
  NOR2X1 U133 ( .A(n79), .B(n85), .Y(\ab[0][4] ) );
  NOR2X1 U134 ( .A(n78), .B(n85), .Y(\ab[0][3] ) );
  NOR2X1 U135 ( .A(n76), .B(n85), .Y(\ab[0][2] ) );
  NOR2X1 U136 ( .A(n74), .B(n85), .Y(\ab[0][1] ) );
  NOR2X1 U137 ( .A(n71), .B(n85), .Y(PRODUCT[0]) );
  INVX2 U99 ( .A(B[0]), .Y(n71) );
  INVX2 U100 ( .A(n49), .Y(n72) );
  INVX2 U101 ( .A(\A1[7] ), .Y(n73) );
  INVX2 U102 ( .A(B[1]), .Y(n74) );
  INVX2 U103 ( .A(n52), .Y(n75) );
  INVX2 U104 ( .A(B[2]), .Y(n76) );
  INVX2 U105 ( .A(n48), .Y(n77) );
  INVX2 U106 ( .A(B[3]), .Y(n78) );
  INVX2 U107 ( .A(B[4]), .Y(n79) );
  INVX2 U108 ( .A(B[5]), .Y(n80) );
  INVX2 U109 ( .A(B[6]), .Y(n81) );
  INVX2 U110 ( .A(B[7]), .Y(n82) );
  INVX2 U111 ( .A(A[2]), .Y(n83) );
  INVX2 U112 ( .A(A[1]), .Y(n84) );
  INVX2 U113 ( .A(A[0]), .Y(n85) );
endmodule


module CannyEdge_DW01_add_39 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_17 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][7] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n61, n62, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n21), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n19), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n18), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n17), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n16), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n15), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(n23), .B(n67), .Y(n3) );
  AND2X2 U3 ( .A(n37), .B(\SUMB[3][2] ), .Y(n4) );
  AND2X2 U4 ( .A(n38), .B(\SUMB[3][3] ), .Y(n5) );
  AND2X2 U5 ( .A(n39), .B(\SUMB[3][4] ), .Y(n6) );
  AND2X2 U6 ( .A(n40), .B(\SUMB[3][5] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[6][1] ), .Y(n8) );
  AND2X2 U8 ( .A(n28), .B(\SUMB[6][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n29), .B(\SUMB[6][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n30), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n32), .B(\SUMB[6][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n41), .B(\CARRYB[2][6] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[4][1] ), .B(n35), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n13), .B(n67), .Y(n22) );
  AND2X2 U22 ( .A(n22), .B(n67), .Y(n23) );
  AND2X2 U23 ( .A(QA), .B(QB), .Y(n24) );
  AND2X2 U24 ( .A(n4), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n5), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n6), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n25), .B(\SUMB[5][2] ), .Y(n28) );
  AND2X2 U28 ( .A(n26), .B(\SUMB[5][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n27), .B(\SUMB[5][4] ), .Y(n30) );
  AND2X2 U30 ( .A(n7), .B(\SUMB[4][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n31), .B(\SUMB[5][5] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][1] ), .B(n8), .Y(n34) );
  AND2X2 U34 ( .A(\SUMB[3][1] ), .B(n33), .Y(n35) );
  AND2X2 U35 ( .A(\SUMB[5][1] ), .B(n14), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n39) );
  AND2X2 U39 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n40) );
  AND2X2 U40 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n67), .Y(n42) );
  AND2X2 U42 ( .A(n67), .B(n3), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n9), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n11), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n12), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n8), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n9), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n10), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n12), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n67), .B(n3), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n24), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U55 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U56 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U57 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U58 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U59 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U60 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U61 ( .A(\SUMB[7][0] ), .B(n67), .Y(\A1[5] ) );
  XOR2X1 U62 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U63 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U64 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U65 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U66 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U67 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U68 ( .A(\SUMB[3][1] ), .B(n33), .Y(\A1[2] ) );
  XOR2X1 U69 ( .A(\SUMB[3][2] ), .B(n37), .Y(\SUMB[4][1] ) );
  XOR2X1 U70 ( .A(\SUMB[3][3] ), .B(n38), .Y(\SUMB[4][2] ) );
  XOR2X1 U71 ( .A(\SUMB[3][4] ), .B(n39), .Y(\SUMB[4][3] ) );
  XOR2X1 U72 ( .A(\SUMB[3][5] ), .B(n40), .Y(\SUMB[4][4] ) );
  XOR2X1 U73 ( .A(\CARRYB[2][6] ), .B(n41), .Y(\SUMB[4][5] ) );
  XOR2X1 U74 ( .A(\SUMB[4][1] ), .B(n35), .Y(\A1[3] ) );
  XOR2X1 U75 ( .A(\SUMB[4][2] ), .B(n4), .Y(\SUMB[5][1] ) );
  XOR2X1 U76 ( .A(\SUMB[4][3] ), .B(n5), .Y(\SUMB[5][2] ) );
  XOR2X1 U77 ( .A(\SUMB[4][4] ), .B(n6), .Y(\SUMB[5][3] ) );
  XOR2X1 U78 ( .A(\SUMB[4][5] ), .B(n7), .Y(\SUMB[5][4] ) );
  XOR2X1 U79 ( .A(n67), .B(n13), .Y(\SUMB[5][5] ) );
  XOR2X1 U80 ( .A(\SUMB[5][1] ), .B(n14), .Y(\A1[4] ) );
  XOR2X1 U81 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U82 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U83 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U84 ( .A(\SUMB[5][5] ), .B(n31), .Y(\SUMB[6][4] ) );
  XOR2X1 U85 ( .A(n67), .B(n22), .Y(\SUMB[6][5] ) );
  XOR2X1 U86 ( .A(\SUMB[6][1] ), .B(n36), .Y(\SUMB[7][0] ) );
  XOR2X1 U87 ( .A(\SUMB[6][2] ), .B(n28), .Y(\SUMB[7][1] ) );
  XOR2X1 U88 ( .A(\SUMB[6][3] ), .B(n29), .Y(\SUMB[7][2] ) );
  XOR2X1 U89 ( .A(\SUMB[6][4] ), .B(n30), .Y(\SUMB[7][3] ) );
  XOR2X1 U90 ( .A(\SUMB[6][5] ), .B(n32), .Y(\SUMB[7][4] ) );
  XOR2X1 U91 ( .A(n67), .B(n23), .Y(\SUMB[7][5] ) );
  XOR2X1 U92 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  NOR2X1 U105 ( .A(n66), .B(n73), .Y(\ab[2][6] ) );
  NOR2X1 U106 ( .A(n66), .B(n72), .Y(\ab[2][5] ) );
  NOR2X1 U107 ( .A(n66), .B(n71), .Y(\ab[2][4] ) );
  NOR2X1 U108 ( .A(n66), .B(n70), .Y(\ab[2][3] ) );
  NOR2X1 U109 ( .A(n66), .B(n69), .Y(\ab[2][2] ) );
  NOR2X1 U110 ( .A(n66), .B(n68), .Y(\ab[2][1] ) );
  NOR2X1 U111 ( .A(n66), .B(n75), .Y(\ab[2][0] ) );
  MUX2X1 U112 ( .B(n61), .A(n62), .S(A[1]), .Y(\ab[1][7] ) );
  NOR2X1 U113 ( .A(n73), .B(n76), .Y(\ab[1][6] ) );
  NOR2X1 U114 ( .A(n72), .B(n76), .Y(\ab[1][5] ) );
  NOR2X1 U115 ( .A(n71), .B(n76), .Y(\ab[1][4] ) );
  NOR2X1 U116 ( .A(n70), .B(n76), .Y(\ab[1][3] ) );
  NOR2X1 U117 ( .A(n69), .B(n76), .Y(\ab[1][2] ) );
  NOR2X1 U118 ( .A(n68), .B(n76), .Y(\ab[1][1] ) );
  NOR2X1 U119 ( .A(n75), .B(n76), .Y(\ab[1][0] ) );
  MUX2X1 U120 ( .B(n61), .A(n62), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U121 ( .A(B[7]), .B(n66), .Y(n62) );
  NOR2X1 U122 ( .A(n73), .B(n74), .Y(\ab[0][6] ) );
  NOR2X1 U123 ( .A(n72), .B(n74), .Y(\ab[0][5] ) );
  NOR2X1 U124 ( .A(n71), .B(n74), .Y(\ab[0][4] ) );
  NOR2X1 U125 ( .A(n70), .B(n74), .Y(\ab[0][3] ) );
  NOR2X1 U126 ( .A(n69), .B(n74), .Y(\ab[0][2] ) );
  NOR2X1 U127 ( .A(n68), .B(n74), .Y(\ab[0][1] ) );
  NAND2X1 U128 ( .A(QA), .B(B[7]), .Y(n61) );
  NOR2X1 U129 ( .A(B[7]), .B(n66), .Y(QB) );
  NOR2X1 U130 ( .A(n75), .B(n74), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_39 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n34, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n66) );
  INVX2 U97 ( .A(n61), .Y(n67) );
  INVX2 U98 ( .A(B[1]), .Y(n68) );
  INVX2 U99 ( .A(B[2]), .Y(n69) );
  INVX2 U100 ( .A(B[3]), .Y(n70) );
  INVX2 U101 ( .A(B[4]), .Y(n71) );
  INVX2 U102 ( .A(B[5]), .Y(n72) );
  INVX2 U103 ( .A(B[6]), .Y(n73) );
  INVX2 U104 ( .A(A[0]), .Y(n74) );
  INVX2 U131 ( .A(B[0]), .Y(n75) );
  INVX2 U132 ( .A(A[1]), .Y(n76) );
endmodule


module CannyEdge_DW01_add_40 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_18 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][7] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n61, n62, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n21), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n19), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n18), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n17), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n16), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n15), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(n23), .B(n67), .Y(n3) );
  AND2X2 U3 ( .A(n36), .B(\SUMB[3][2] ), .Y(n4) );
  AND2X2 U4 ( .A(n37), .B(\SUMB[3][3] ), .Y(n5) );
  AND2X2 U5 ( .A(n38), .B(\SUMB[3][4] ), .Y(n6) );
  AND2X2 U6 ( .A(n39), .B(\SUMB[3][5] ), .Y(n7) );
  AND2X2 U7 ( .A(n35), .B(\SUMB[6][1] ), .Y(n8) );
  AND2X2 U8 ( .A(n27), .B(\SUMB[6][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n28), .B(\SUMB[6][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n29), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n31), .B(\SUMB[6][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n40), .B(\CARRYB[2][6] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[4][1] ), .B(n34), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n13), .B(n67), .Y(n22) );
  AND2X2 U22 ( .A(n22), .B(n67), .Y(n23) );
  AND2X2 U23 ( .A(n4), .B(\SUMB[4][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n5), .B(\SUMB[4][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n6), .B(\SUMB[4][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n24), .B(\SUMB[5][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n25), .B(\SUMB[5][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n26), .B(\SUMB[5][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n7), .B(\SUMB[4][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n30), .B(\SUMB[5][5] ), .Y(n31) );
  AND2X2 U31 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][1] ), .B(n8), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[3][1] ), .B(n32), .Y(n34) );
  AND2X2 U34 ( .A(\SUMB[5][1] ), .B(n14), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n39) );
  AND2X2 U39 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n40) );
  AND2X2 U40 ( .A(QA), .B(QB), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n67), .Y(n42) );
  AND2X2 U42 ( .A(n67), .B(n3), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n9), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n11), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n12), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n8), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n9), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n10), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n12), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n67), .B(n3), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n41), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U55 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U56 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U57 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U58 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U59 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U60 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U61 ( .A(\SUMB[7][0] ), .B(n67), .Y(\A1[5] ) );
  XOR2X1 U62 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U63 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U64 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U65 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U66 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U67 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U68 ( .A(\SUMB[3][1] ), .B(n32), .Y(\A1[2] ) );
  XOR2X1 U69 ( .A(\SUMB[3][2] ), .B(n36), .Y(\SUMB[4][1] ) );
  XOR2X1 U70 ( .A(\SUMB[3][3] ), .B(n37), .Y(\SUMB[4][2] ) );
  XOR2X1 U71 ( .A(\SUMB[3][4] ), .B(n38), .Y(\SUMB[4][3] ) );
  XOR2X1 U72 ( .A(\SUMB[3][5] ), .B(n39), .Y(\SUMB[4][4] ) );
  XOR2X1 U73 ( .A(\CARRYB[2][6] ), .B(n40), .Y(\SUMB[4][5] ) );
  XOR2X1 U74 ( .A(\SUMB[4][1] ), .B(n34), .Y(\A1[3] ) );
  XOR2X1 U75 ( .A(\SUMB[4][2] ), .B(n4), .Y(\SUMB[5][1] ) );
  XOR2X1 U76 ( .A(\SUMB[4][3] ), .B(n5), .Y(\SUMB[5][2] ) );
  XOR2X1 U77 ( .A(\SUMB[4][4] ), .B(n6), .Y(\SUMB[5][3] ) );
  XOR2X1 U78 ( .A(\SUMB[4][5] ), .B(n7), .Y(\SUMB[5][4] ) );
  XOR2X1 U79 ( .A(n67), .B(n13), .Y(\SUMB[5][5] ) );
  XOR2X1 U80 ( .A(\SUMB[5][1] ), .B(n14), .Y(\A1[4] ) );
  XOR2X1 U81 ( .A(\SUMB[5][2] ), .B(n24), .Y(\SUMB[6][1] ) );
  XOR2X1 U82 ( .A(\SUMB[5][3] ), .B(n25), .Y(\SUMB[6][2] ) );
  XOR2X1 U83 ( .A(\SUMB[5][4] ), .B(n26), .Y(\SUMB[6][3] ) );
  XOR2X1 U84 ( .A(\SUMB[5][5] ), .B(n30), .Y(\SUMB[6][4] ) );
  XOR2X1 U85 ( .A(n67), .B(n22), .Y(\SUMB[6][5] ) );
  XOR2X1 U86 ( .A(\SUMB[6][1] ), .B(n35), .Y(\SUMB[7][0] ) );
  XOR2X1 U87 ( .A(\SUMB[6][2] ), .B(n27), .Y(\SUMB[7][1] ) );
  XOR2X1 U88 ( .A(\SUMB[6][3] ), .B(n28), .Y(\SUMB[7][2] ) );
  XOR2X1 U89 ( .A(\SUMB[6][4] ), .B(n29), .Y(\SUMB[7][3] ) );
  XOR2X1 U90 ( .A(\SUMB[6][5] ), .B(n31), .Y(\SUMB[7][4] ) );
  XOR2X1 U91 ( .A(n67), .B(n23), .Y(\SUMB[7][5] ) );
  XOR2X1 U92 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  NOR2X1 U105 ( .A(n66), .B(n73), .Y(\ab[2][6] ) );
  NOR2X1 U106 ( .A(n66), .B(n72), .Y(\ab[2][5] ) );
  NOR2X1 U107 ( .A(n66), .B(n71), .Y(\ab[2][4] ) );
  NOR2X1 U108 ( .A(n66), .B(n70), .Y(\ab[2][3] ) );
  NOR2X1 U109 ( .A(n66), .B(n69), .Y(\ab[2][2] ) );
  NOR2X1 U110 ( .A(n66), .B(n68), .Y(\ab[2][1] ) );
  NOR2X1 U111 ( .A(n66), .B(n75), .Y(\ab[2][0] ) );
  MUX2X1 U112 ( .B(n61), .A(n62), .S(A[1]), .Y(\ab[1][7] ) );
  NOR2X1 U113 ( .A(n73), .B(n76), .Y(\ab[1][6] ) );
  NOR2X1 U114 ( .A(n72), .B(n76), .Y(\ab[1][5] ) );
  NOR2X1 U115 ( .A(n71), .B(n76), .Y(\ab[1][4] ) );
  NOR2X1 U116 ( .A(n70), .B(n76), .Y(\ab[1][3] ) );
  NOR2X1 U117 ( .A(n69), .B(n76), .Y(\ab[1][2] ) );
  NOR2X1 U118 ( .A(n68), .B(n76), .Y(\ab[1][1] ) );
  NOR2X1 U119 ( .A(n75), .B(n76), .Y(\ab[1][0] ) );
  MUX2X1 U120 ( .B(n61), .A(n62), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U121 ( .A(B[7]), .B(n66), .Y(n62) );
  NOR2X1 U122 ( .A(n73), .B(n74), .Y(\ab[0][6] ) );
  NOR2X1 U123 ( .A(n72), .B(n74), .Y(\ab[0][5] ) );
  NOR2X1 U124 ( .A(n71), .B(n74), .Y(\ab[0][4] ) );
  NOR2X1 U125 ( .A(n70), .B(n74), .Y(\ab[0][3] ) );
  NOR2X1 U126 ( .A(n69), .B(n74), .Y(\ab[0][2] ) );
  NOR2X1 U127 ( .A(n68), .B(n74), .Y(\ab[0][1] ) );
  NAND2X1 U128 ( .A(QA), .B(B[7]), .Y(n61) );
  NOR2X1 U129 ( .A(B[7]), .B(n66), .Y(QB) );
  NOR2X1 U130 ( .A(n75), .B(n74), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_40 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n33, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n66) );
  INVX2 U97 ( .A(n61), .Y(n67) );
  INVX2 U98 ( .A(B[1]), .Y(n68) );
  INVX2 U99 ( .A(B[2]), .Y(n69) );
  INVX2 U100 ( .A(B[3]), .Y(n70) );
  INVX2 U101 ( .A(B[4]), .Y(n71) );
  INVX2 U102 ( .A(B[5]), .Y(n72) );
  INVX2 U103 ( .A(B[6]), .Y(n73) );
  INVX2 U104 ( .A(A[0]), .Y(n74) );
  INVX2 U131 ( .A(B[0]), .Y(n75) );
  INVX2 U132 ( .A(A[1]), .Y(n76) );
endmodule


module CannyEdge_DW01_cmp2_3 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174;

  AND2X2 U1 ( .A(n130), .B(n60), .Y(n1) );
  MUX2X1 U59 ( .B(n1), .A(TC), .S(A[31]), .Y(GE_GT) );
  AOI21X1 U60 ( .A(A[29]), .B(n173), .C(n61), .Y(n60) );
  AOI21X1 U61 ( .A(B[29]), .B(n131), .C(n62), .Y(n61) );
  OAI21X1 U62 ( .A(A[28]), .B(n172), .C(n63), .Y(n62) );
  OAI21X1 U63 ( .A(B[28]), .B(n132), .C(n64), .Y(n63) );
  AOI21X1 U64 ( .A(A[27]), .B(n171), .C(n65), .Y(n64) );
  AOI21X1 U65 ( .A(B[27]), .B(n133), .C(n66), .Y(n65) );
  OAI21X1 U66 ( .A(A[26]), .B(n170), .C(n67), .Y(n66) );
  OAI21X1 U67 ( .A(B[26]), .B(n134), .C(n68), .Y(n67) );
  AOI21X1 U68 ( .A(A[25]), .B(n169), .C(n69), .Y(n68) );
  AOI21X1 U69 ( .A(B[25]), .B(n135), .C(n70), .Y(n69) );
  OAI21X1 U70 ( .A(A[24]), .B(n168), .C(n71), .Y(n70) );
  OAI21X1 U71 ( .A(B[24]), .B(n136), .C(n72), .Y(n71) );
  AOI21X1 U72 ( .A(A[23]), .B(n167), .C(n73), .Y(n72) );
  AOI21X1 U73 ( .A(B[23]), .B(n137), .C(n74), .Y(n73) );
  OAI21X1 U74 ( .A(A[22]), .B(n166), .C(n75), .Y(n74) );
  OAI21X1 U75 ( .A(B[22]), .B(n138), .C(n76), .Y(n75) );
  AOI21X1 U76 ( .A(A[21]), .B(n165), .C(n77), .Y(n76) );
  AOI21X1 U77 ( .A(B[21]), .B(n139), .C(n78), .Y(n77) );
  OAI21X1 U78 ( .A(A[20]), .B(n164), .C(n79), .Y(n78) );
  OAI21X1 U79 ( .A(B[20]), .B(n140), .C(n80), .Y(n79) );
  AOI21X1 U80 ( .A(A[19]), .B(n163), .C(n81), .Y(n80) );
  AOI21X1 U81 ( .A(B[19]), .B(n141), .C(n82), .Y(n81) );
  OAI21X1 U82 ( .A(A[18]), .B(n162), .C(n83), .Y(n82) );
  OAI21X1 U83 ( .A(B[18]), .B(n142), .C(n84), .Y(n83) );
  AOI21X1 U84 ( .A(A[17]), .B(n161), .C(n85), .Y(n84) );
  AOI21X1 U85 ( .A(B[17]), .B(n143), .C(n86), .Y(n85) );
  OAI21X1 U86 ( .A(A[16]), .B(n160), .C(n87), .Y(n86) );
  OAI21X1 U87 ( .A(B[16]), .B(n144), .C(n88), .Y(n87) );
  AOI21X1 U88 ( .A(A[15]), .B(n159), .C(n89), .Y(n88) );
  AOI21X1 U89 ( .A(B[15]), .B(n145), .C(n90), .Y(n89) );
  OAI21X1 U90 ( .A(A[14]), .B(n158), .C(n91), .Y(n90) );
  OAI21X1 U91 ( .A(B[14]), .B(n146), .C(n92), .Y(n91) );
  AOI21X1 U92 ( .A(A[13]), .B(n157), .C(n93), .Y(n92) );
  AOI21X1 U93 ( .A(B[13]), .B(n147), .C(n94), .Y(n93) );
  OAI21X1 U94 ( .A(A[12]), .B(n156), .C(n95), .Y(n94) );
  OAI21X1 U95 ( .A(B[12]), .B(n148), .C(n96), .Y(n95) );
  AOI21X1 U96 ( .A(A[11]), .B(n155), .C(n97), .Y(n96) );
  AOI21X1 U97 ( .A(B[11]), .B(n149), .C(n98), .Y(n97) );
  OAI21X1 U98 ( .A(A[10]), .B(n154), .C(n99), .Y(n98) );
  OAI21X1 U99 ( .A(B[9]), .B(n128), .C(n100), .Y(n99) );
  AOI21X1 U100 ( .A(A[10]), .B(n154), .C(n101), .Y(n100) );
  AOI21X1 U101 ( .A(B[9]), .B(n128), .C(n102), .Y(n101) );
  OAI21X1 U102 ( .A(A[8]), .B(n174), .C(n103), .Y(n102) );
  OAI21X1 U103 ( .A(B[8]), .B(n129), .C(n104), .Y(n103) );
  AOI21X1 U104 ( .A(A[7]), .B(n118), .C(n105), .Y(n104) );
  AOI21X1 U105 ( .A(B[7]), .B(n150), .C(n106), .Y(n105) );
  OAI21X1 U106 ( .A(A[6]), .B(n119), .C(n107), .Y(n106) );
  OAI21X1 U107 ( .A(B[6]), .B(n151), .C(n108), .Y(n107) );
  AOI21X1 U108 ( .A(A[5]), .B(n120), .C(n109), .Y(n108) );
  AOI21X1 U109 ( .A(B[5]), .B(n152), .C(n110), .Y(n109) );
  OAI21X1 U110 ( .A(A[4]), .B(n121), .C(n111), .Y(n110) );
  OAI21X1 U111 ( .A(B[4]), .B(n153), .C(n112), .Y(n111) );
  AOI21X1 U112 ( .A(A[3]), .B(n122), .C(n113), .Y(n112) );
  AOI21X1 U113 ( .A(B[3]), .B(n127), .C(n114), .Y(n113) );
  OAI21X1 U114 ( .A(A[2]), .B(n123), .C(n115), .Y(n114) );
  OAI21X1 U115 ( .A(B[2]), .B(n126), .C(n116), .Y(n115) );
  AOI22X1 U116 ( .A(n117), .B(A[0]), .C(A[1]), .D(n124), .Y(n116) );
  AOI21X1 U117 ( .A(B[1]), .B(n125), .C(B[0]), .Y(n117) );
  INVX2 U2 ( .A(B[7]), .Y(n118) );
  INVX2 U3 ( .A(B[6]), .Y(n119) );
  INVX2 U4 ( .A(B[5]), .Y(n120) );
  INVX2 U5 ( .A(B[4]), .Y(n121) );
  INVX2 U6 ( .A(B[3]), .Y(n122) );
  INVX2 U7 ( .A(B[2]), .Y(n123) );
  INVX2 U8 ( .A(B[1]), .Y(n124) );
  INVX2 U9 ( .A(A[1]), .Y(n125) );
  INVX2 U10 ( .A(A[2]), .Y(n126) );
  INVX2 U11 ( .A(A[3]), .Y(n127) );
  INVX2 U12 ( .A(A[9]), .Y(n128) );
  INVX2 U13 ( .A(A[8]), .Y(n129) );
  INVX2 U14 ( .A(A[30]), .Y(n130) );
  INVX2 U15 ( .A(A[29]), .Y(n131) );
  INVX2 U16 ( .A(A[28]), .Y(n132) );
  INVX2 U17 ( .A(A[27]), .Y(n133) );
  INVX2 U18 ( .A(A[26]), .Y(n134) );
  INVX2 U19 ( .A(A[25]), .Y(n135) );
  INVX2 U20 ( .A(A[24]), .Y(n136) );
  INVX2 U21 ( .A(A[23]), .Y(n137) );
  INVX2 U22 ( .A(A[22]), .Y(n138) );
  INVX2 U23 ( .A(A[21]), .Y(n139) );
  INVX2 U24 ( .A(A[20]), .Y(n140) );
  INVX2 U25 ( .A(A[19]), .Y(n141) );
  INVX2 U26 ( .A(A[18]), .Y(n142) );
  INVX2 U27 ( .A(A[17]), .Y(n143) );
  INVX2 U28 ( .A(A[16]), .Y(n144) );
  INVX2 U29 ( .A(A[15]), .Y(n145) );
  INVX2 U30 ( .A(A[14]), .Y(n146) );
  INVX2 U31 ( .A(A[13]), .Y(n147) );
  INVX2 U32 ( .A(A[12]), .Y(n148) );
  INVX2 U33 ( .A(A[11]), .Y(n149) );
  INVX2 U34 ( .A(A[7]), .Y(n150) );
  INVX2 U35 ( .A(A[6]), .Y(n151) );
  INVX2 U36 ( .A(A[5]), .Y(n152) );
  INVX2 U37 ( .A(A[4]), .Y(n153) );
  INVX2 U38 ( .A(B[10]), .Y(n154) );
  INVX2 U39 ( .A(B[11]), .Y(n155) );
  INVX2 U40 ( .A(B[12]), .Y(n156) );
  INVX2 U41 ( .A(B[13]), .Y(n157) );
  INVX2 U42 ( .A(B[14]), .Y(n158) );
  INVX2 U43 ( .A(B[15]), .Y(n159) );
  INVX2 U44 ( .A(B[16]), .Y(n160) );
  INVX2 U45 ( .A(B[17]), .Y(n161) );
  INVX2 U46 ( .A(B[18]), .Y(n162) );
  INVX2 U47 ( .A(B[19]), .Y(n163) );
  INVX2 U48 ( .A(B[20]), .Y(n164) );
  INVX2 U49 ( .A(B[21]), .Y(n165) );
  INVX2 U50 ( .A(B[22]), .Y(n166) );
  INVX2 U51 ( .A(B[23]), .Y(n167) );
  INVX2 U52 ( .A(B[24]), .Y(n168) );
  INVX2 U53 ( .A(B[25]), .Y(n169) );
  INVX2 U54 ( .A(B[26]), .Y(n170) );
  INVX2 U55 ( .A(B[27]), .Y(n171) );
  INVX2 U56 ( .A(B[28]), .Y(n172) );
  INVX2 U57 ( .A(B[29]), .Y(n173) );
  INVX2 U58 ( .A(B[8]), .Y(n174) );
endmodule


module CannyEdge_DW01_add_41 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U31 ( .A(n30), .B(n31), .Y(SUM[9]) );
  NOR2X1 U32 ( .A(n127), .B(n32), .Y(n31) );
  XOR2X1 U33 ( .A(n34), .B(n131), .Y(SUM[8]) );
  NAND2X1 U34 ( .A(n130), .B(n35), .Y(n34) );
  XOR2X1 U35 ( .A(n37), .B(n38), .Y(SUM[7]) );
  XOR2X1 U36 ( .A(n132), .B(B[7]), .Y(n38) );
  OAI21X1 U37 ( .A(B[6]), .B(A[6]), .C(n37), .Y(n39) );
  XOR2X1 U38 ( .A(n40), .B(n41), .Y(SUM[29]) );
  XOR2X1 U39 ( .A(B[29]), .B(A[29]), .Y(n41) );
  OAI21X1 U40 ( .A(n42), .B(n43), .C(n44), .Y(n40) );
  XOR2X1 U41 ( .A(n45), .B(n43), .Y(SUM[28]) );
  AOI21X1 U42 ( .A(n148), .B(n46), .C(n47), .Y(n43) );
  NAND2X1 U43 ( .A(n149), .B(n44), .Y(n45) );
  NAND2X1 U44 ( .A(B[28]), .B(A[28]), .Y(n44) );
  NOR2X1 U45 ( .A(B[28]), .B(A[28]), .Y(n42) );
  XOR2X1 U46 ( .A(n46), .B(n49), .Y(SUM[27]) );
  NOR2X1 U47 ( .A(n47), .B(n48), .Y(n49) );
  NOR2X1 U48 ( .A(B[27]), .B(A[27]), .Y(n48) );
  AND2X1 U49 ( .A(B[27]), .B(A[27]), .Y(n47) );
  OAI21X1 U50 ( .A(n50), .B(n51), .C(n52), .Y(n46) );
  XOR2X1 U51 ( .A(n53), .B(n51), .Y(SUM[26]) );
  AOI21X1 U52 ( .A(n146), .B(n54), .C(n55), .Y(n51) );
  NAND2X1 U53 ( .A(n147), .B(n52), .Y(n53) );
  NAND2X1 U54 ( .A(B[26]), .B(A[26]), .Y(n52) );
  NOR2X1 U55 ( .A(B[26]), .B(A[26]), .Y(n50) );
  XOR2X1 U56 ( .A(n54), .B(n57), .Y(SUM[25]) );
  NOR2X1 U57 ( .A(n55), .B(n56), .Y(n57) );
  NOR2X1 U58 ( .A(B[25]), .B(A[25]), .Y(n56) );
  AND2X1 U59 ( .A(B[25]), .B(A[25]), .Y(n55) );
  OAI21X1 U60 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  XOR2X1 U61 ( .A(n61), .B(n59), .Y(SUM[24]) );
  AOI21X1 U62 ( .A(n144), .B(n62), .C(n63), .Y(n59) );
  NAND2X1 U63 ( .A(n145), .B(n60), .Y(n61) );
  NAND2X1 U64 ( .A(B[24]), .B(A[24]), .Y(n60) );
  NOR2X1 U65 ( .A(B[24]), .B(A[24]), .Y(n58) );
  XOR2X1 U66 ( .A(n62), .B(n65), .Y(SUM[23]) );
  NOR2X1 U67 ( .A(n63), .B(n64), .Y(n65) );
  NOR2X1 U68 ( .A(B[23]), .B(A[23]), .Y(n64) );
  AND2X1 U69 ( .A(B[23]), .B(A[23]), .Y(n63) );
  OAI21X1 U70 ( .A(n66), .B(n67), .C(n68), .Y(n62) );
  XOR2X1 U71 ( .A(n69), .B(n67), .Y(SUM[22]) );
  AOI21X1 U72 ( .A(n142), .B(n70), .C(n71), .Y(n67) );
  NAND2X1 U73 ( .A(n143), .B(n68), .Y(n69) );
  NAND2X1 U74 ( .A(B[22]), .B(A[22]), .Y(n68) );
  NOR2X1 U75 ( .A(B[22]), .B(A[22]), .Y(n66) );
  XOR2X1 U76 ( .A(n70), .B(n73), .Y(SUM[21]) );
  NOR2X1 U77 ( .A(n71), .B(n72), .Y(n73) );
  NOR2X1 U78 ( .A(B[21]), .B(A[21]), .Y(n72) );
  AND2X1 U79 ( .A(B[21]), .B(A[21]), .Y(n71) );
  OAI21X1 U80 ( .A(n74), .B(n75), .C(n76), .Y(n70) );
  XOR2X1 U81 ( .A(n77), .B(n75), .Y(SUM[20]) );
  AOI21X1 U82 ( .A(n140), .B(n78), .C(n79), .Y(n75) );
  NAND2X1 U83 ( .A(n141), .B(n76), .Y(n77) );
  NAND2X1 U84 ( .A(B[20]), .B(A[20]), .Y(n76) );
  NOR2X1 U85 ( .A(B[20]), .B(A[20]), .Y(n74) );
  XOR2X1 U86 ( .A(n78), .B(n81), .Y(SUM[19]) );
  NOR2X1 U87 ( .A(n79), .B(n80), .Y(n81) );
  NOR2X1 U88 ( .A(B[19]), .B(A[19]), .Y(n80) );
  AND2X1 U89 ( .A(B[19]), .B(A[19]), .Y(n79) );
  OAI21X1 U90 ( .A(n82), .B(n83), .C(n84), .Y(n78) );
  XOR2X1 U91 ( .A(n85), .B(n83), .Y(SUM[18]) );
  AOI21X1 U92 ( .A(n136), .B(n86), .C(n87), .Y(n83) );
  NAND2X1 U93 ( .A(n139), .B(n84), .Y(n85) );
  NAND2X1 U94 ( .A(B[18]), .B(A[18]), .Y(n84) );
  NOR2X1 U95 ( .A(B[18]), .B(A[18]), .Y(n82) );
  XOR2X1 U96 ( .A(n86), .B(n89), .Y(SUM[17]) );
  NOR2X1 U97 ( .A(n87), .B(n88), .Y(n89) );
  NOR2X1 U98 ( .A(B[17]), .B(A[17]), .Y(n88) );
  AND2X1 U99 ( .A(B[17]), .B(A[17]), .Y(n87) );
  OAI21X1 U100 ( .A(n90), .B(n91), .C(n92), .Y(n86) );
  XOR2X1 U101 ( .A(n93), .B(n91), .Y(SUM[16]) );
  AOI21X1 U102 ( .A(n138), .B(n94), .C(n95), .Y(n91) );
  NAND2X1 U103 ( .A(n137), .B(n92), .Y(n93) );
  NAND2X1 U104 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NOR2X1 U105 ( .A(B[16]), .B(A[16]), .Y(n90) );
  XOR2X1 U106 ( .A(n94), .B(n97), .Y(SUM[15]) );
  NOR2X1 U107 ( .A(n95), .B(n96), .Y(n97) );
  NOR2X1 U108 ( .A(B[15]), .B(A[15]), .Y(n96) );
  AND2X1 U109 ( .A(B[15]), .B(A[15]), .Y(n95) );
  OAI21X1 U110 ( .A(n98), .B(n99), .C(n100), .Y(n94) );
  XOR2X1 U111 ( .A(n101), .B(n99), .Y(SUM[14]) );
  AOI21X1 U112 ( .A(n121), .B(n102), .C(n103), .Y(n99) );
  NAND2X1 U113 ( .A(n135), .B(n100), .Y(n101) );
  NAND2X1 U114 ( .A(B[14]), .B(A[14]), .Y(n100) );
  NOR2X1 U115 ( .A(B[14]), .B(A[14]), .Y(n98) );
  XOR2X1 U116 ( .A(n102), .B(n105), .Y(SUM[13]) );
  NOR2X1 U117 ( .A(n103), .B(n104), .Y(n105) );
  NOR2X1 U118 ( .A(B[13]), .B(A[13]), .Y(n104) );
  AND2X1 U119 ( .A(B[13]), .B(A[13]), .Y(n103) );
  OAI21X1 U120 ( .A(n106), .B(n123), .C(n107), .Y(n102) );
  XOR2X1 U121 ( .A(n108), .B(n123), .Y(SUM[12]) );
  OAI21X1 U122 ( .A(n110), .B(n111), .C(n112), .Y(n109) );
  AOI21X1 U123 ( .A(n113), .B(n126), .C(n125), .Y(n111) );
  NAND2X1 U124 ( .A(n122), .B(n107), .Y(n108) );
  NAND2X1 U125 ( .A(B[12]), .B(A[12]), .Y(n107) );
  NOR2X1 U126 ( .A(B[12]), .B(A[12]), .Y(n106) );
  XOR2X1 U127 ( .A(n115), .B(n116), .Y(SUM[11]) );
  NOR2X1 U128 ( .A(n124), .B(n110), .Y(n116) );
  NOR2X1 U129 ( .A(B[11]), .B(A[11]), .Y(n110) );
  NAND2X1 U130 ( .A(B[11]), .B(A[11]), .Y(n112) );
  OAI21X1 U131 ( .A(n117), .B(n128), .C(n114), .Y(n115) );
  XOR2X1 U132 ( .A(n118), .B(n128), .Y(SUM[10]) );
  OAI21X1 U133 ( .A(n129), .B(n32), .C(n33), .Y(n113) );
  NAND2X1 U134 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NOR2X1 U135 ( .A(B[9]), .B(A[9]), .Y(n32) );
  OAI21X1 U136 ( .A(n36), .B(n131), .C(n35), .Y(n30) );
  NAND2X1 U137 ( .A(B[8]), .B(A[8]), .Y(n35) );
  OAI21X1 U138 ( .A(n37), .B(n132), .C(n120), .Y(n119) );
  OAI21X1 U139 ( .A(n134), .B(A[7]), .C(B[7]), .Y(n120) );
  NAND2X1 U140 ( .A(B[6]), .B(A[6]), .Y(n37) );
  NOR2X1 U141 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NAND2X1 U142 ( .A(n126), .B(n114), .Y(n118) );
  NAND2X1 U143 ( .A(B[10]), .B(A[10]), .Y(n114) );
  NOR2X1 U144 ( .A(B[10]), .B(A[10]), .Y(n117) );
  INVX2 U2 ( .A(n104), .Y(n121) );
  INVX2 U3 ( .A(n106), .Y(n122) );
  INVX2 U4 ( .A(n109), .Y(n123) );
  INVX2 U5 ( .A(n112), .Y(n124) );
  INVX2 U6 ( .A(n114), .Y(n125) );
  INVX2 U7 ( .A(n117), .Y(n126) );
  INVX2 U8 ( .A(n33), .Y(n127) );
  INVX2 U9 ( .A(n113), .Y(n128) );
  INVX2 U10 ( .A(n30), .Y(n129) );
  INVX2 U11 ( .A(n36), .Y(n130) );
  INVX2 U12 ( .A(n119), .Y(n131) );
  INVX2 U13 ( .A(A[7]), .Y(n132) );
  INVX2 U14 ( .A(n39), .Y(SUM[6]) );
  INVX2 U15 ( .A(n37), .Y(n134) );
  INVX2 U16 ( .A(n98), .Y(n135) );
  INVX2 U17 ( .A(n88), .Y(n136) );
  INVX2 U18 ( .A(n90), .Y(n137) );
  INVX2 U19 ( .A(n96), .Y(n138) );
  INVX2 U20 ( .A(n82), .Y(n139) );
  INVX2 U21 ( .A(n80), .Y(n140) );
  INVX2 U22 ( .A(n74), .Y(n141) );
  INVX2 U23 ( .A(n72), .Y(n142) );
  INVX2 U24 ( .A(n66), .Y(n143) );
  INVX2 U25 ( .A(n64), .Y(n144) );
  INVX2 U26 ( .A(n58), .Y(n145) );
  INVX2 U27 ( .A(n56), .Y(n146) );
  INVX2 U28 ( .A(n50), .Y(n147) );
  INVX2 U29 ( .A(n48), .Y(n148) );
  INVX2 U30 ( .A(n42), .Y(n149) );
endmodule


module CannyEdge_DW02_mult_19 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] , \ab[7][27] ,
         \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][31] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][31] , \ab[3][30] ,
         \ab[3][29] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] , \ab[2][27] ,
         \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][31] ,
         \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] ,
         \ab[0][25] , \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] ,
         \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] ,
         \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] ,
         \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] ,
         \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] ,
         \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[30] , n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n110, n111, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S14_31_0 ( .A(n152), .B(\CARRYB[7][23] ), .C(\SUMB[7][24] ), .YC(
        \A2[30] ), .YS(\A1[29] ) );
  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S4_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S4_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S4_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S4_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  FAX1 S4_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S4_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S4_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S4_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  FAX1 S4_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S4_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S4_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S4_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  FAX1 S4_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S4_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S4_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S4_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  FAX1 S4_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S4_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S4_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S4_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  FAX1 S4_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S4_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S5_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .C(\ab[6][31] ), .YC(
        \CARRYB[7][30] ), .YS(\SUMB[7][30] ) );
  FAX1 S14_31 ( .A(QA), .B(QB), .C(\ab[7][31] ), .YC(\CARRYB[7][31] ), .YS(
        \SUMB[7][31] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  FAX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  FAX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  FAX1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  FAX1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  FAX1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .C(\ab[5][31] ), .YC(
        \CARRYB[6][30] ), .YS(\SUMB[6][30] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .C(\ab[4][31] ), .YC(
        \CARRYB[5][30] ), .YS(\SUMB[5][30] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .C(\ab[3][31] ), .YC(
        \CARRYB[4][30] ), .YS(\SUMB[4][30] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .C(\ab[2][31] ), .YC(
        \CARRYB[3][30] ), .YS(\SUMB[3][30] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n42), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n41), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n40), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n39), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n38), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n37), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n36), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n35), .C(\SUMB[1][8] ), .YC(\CARRYB[2][7] ), 
        .YS(\SUMB[2][7] ) );
  FAX1 S2_2_8 ( .A(\ab[2][8] ), .B(n34), .C(\SUMB[1][9] ), .YC(\CARRYB[2][8] ), 
        .YS(\SUMB[2][8] ) );
  FAX1 S2_2_9 ( .A(\ab[2][9] ), .B(n33), .C(\SUMB[1][10] ), .YC(\CARRYB[2][9] ), .YS(\SUMB[2][9] ) );
  FAX1 S2_2_10 ( .A(\ab[2][10] ), .B(n32), .C(\SUMB[1][11] ), .YC(
        \CARRYB[2][10] ), .YS(\SUMB[2][10] ) );
  FAX1 S2_2_11 ( .A(\ab[2][11] ), .B(n31), .C(\SUMB[1][12] ), .YC(
        \CARRYB[2][11] ), .YS(\SUMB[2][11] ) );
  FAX1 S2_2_12 ( .A(\ab[2][12] ), .B(n30), .C(\SUMB[1][13] ), .YC(
        \CARRYB[2][12] ), .YS(\SUMB[2][12] ) );
  FAX1 S2_2_13 ( .A(\ab[2][13] ), .B(n29), .C(\SUMB[1][14] ), .YC(
        \CARRYB[2][13] ), .YS(\SUMB[2][13] ) );
  FAX1 S2_2_14 ( .A(\ab[2][14] ), .B(n28), .C(\SUMB[1][15] ), .YC(
        \CARRYB[2][14] ), .YS(\SUMB[2][14] ) );
  FAX1 S2_2_15 ( .A(\ab[2][15] ), .B(n27), .C(\SUMB[1][16] ), .YC(
        \CARRYB[2][15] ), .YS(\SUMB[2][15] ) );
  FAX1 S2_2_16 ( .A(\ab[2][16] ), .B(n26), .C(\SUMB[1][17] ), .YC(
        \CARRYB[2][16] ), .YS(\SUMB[2][16] ) );
  FAX1 S2_2_17 ( .A(\ab[2][17] ), .B(n25), .C(\SUMB[1][18] ), .YC(
        \CARRYB[2][17] ), .YS(\SUMB[2][17] ) );
  FAX1 S2_2_18 ( .A(\ab[2][18] ), .B(n24), .C(\SUMB[1][19] ), .YC(
        \CARRYB[2][18] ), .YS(\SUMB[2][18] ) );
  FAX1 S2_2_19 ( .A(\ab[2][19] ), .B(n23), .C(\SUMB[1][20] ), .YC(
        \CARRYB[2][19] ), .YS(\SUMB[2][19] ) );
  FAX1 S2_2_20 ( .A(\ab[2][20] ), .B(n22), .C(\SUMB[1][21] ), .YC(
        \CARRYB[2][20] ), .YS(\SUMB[2][20] ) );
  FAX1 S2_2_21 ( .A(\ab[2][21] ), .B(n21), .C(\SUMB[1][22] ), .YC(
        \CARRYB[2][21] ), .YS(\SUMB[2][21] ) );
  FAX1 S2_2_22 ( .A(\ab[2][22] ), .B(n20), .C(\SUMB[1][23] ), .YC(
        \CARRYB[2][22] ), .YS(\SUMB[2][22] ) );
  FAX1 S2_2_23 ( .A(\ab[2][23] ), .B(n19), .C(\SUMB[1][24] ), .YC(
        \CARRYB[2][23] ), .YS(\SUMB[2][23] ) );
  FAX1 S2_2_24 ( .A(\ab[2][24] ), .B(n18), .C(\SUMB[1][25] ), .YC(
        \CARRYB[2][24] ), .YS(\SUMB[2][24] ) );
  FAX1 S2_2_25 ( .A(\ab[2][25] ), .B(n17), .C(\SUMB[1][26] ), .YC(
        \CARRYB[2][25] ), .YS(\SUMB[2][25] ) );
  FAX1 S2_2_26 ( .A(\ab[2][26] ), .B(n16), .C(\SUMB[1][27] ), .YC(
        \CARRYB[2][26] ), .YS(\SUMB[2][26] ) );
  FAX1 S2_2_27 ( .A(\ab[2][27] ), .B(n15), .C(\SUMB[1][28] ), .YC(
        \CARRYB[2][27] ), .YS(\SUMB[2][27] ) );
  FAX1 S2_2_28 ( .A(\ab[2][28] ), .B(n14), .C(\SUMB[1][29] ), .YC(
        \CARRYB[2][28] ), .YS(\SUMB[2][28] ) );
  FAX1 S2_2_29 ( .A(\ab[2][29] ), .B(n13), .C(\SUMB[1][30] ), .YC(
        \CARRYB[2][29] ), .YS(\SUMB[2][29] ) );
  FAX1 S3_2_30 ( .A(\ab[2][30] ), .B(n12), .C(\ab[1][31] ), .YC(
        \CARRYB[2][30] ), .YS(\SUMB[2][30] ) );
  AND2X2 U2 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(n3) );
  AND2X2 U3 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(n4) );
  AND2X2 U4 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(n5) );
  AND2X2 U5 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(n6) );
  AND2X2 U6 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(n7) );
  AND2X2 U7 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(n8) );
  AND2X2 U8 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(n9) );
  AND2X2 U9 ( .A(TC), .B(A[7]), .Y(n10) );
  AND2X2 U10 ( .A(A[7]), .B(n155), .Y(n11) );
  AND2X2 U11 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Y(n12) );
  AND2X2 U12 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Y(n13) );
  AND2X2 U13 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Y(n24) );
  AND2X2 U24 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Y(n25) );
  AND2X2 U25 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Y(n26) );
  AND2X2 U26 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Y(n27) );
  AND2X2 U27 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n28) );
  AND2X2 U28 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n29) );
  AND2X2 U29 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n30) );
  AND2X2 U30 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Y(n31) );
  AND2X2 U31 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n36) );
  AND2X2 U36 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n37) );
  AND2X2 U37 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n38) );
  AND2X2 U38 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n39) );
  AND2X2 U39 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n40) );
  AND2X2 U40 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n41) );
  AND2X2 U41 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n42) );
  AND2X2 U42 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][0] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(n53) );
  AND2X2 U53 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(n54) );
  AND2X2 U54 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(n55) );
  AND2X2 U55 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(n56) );
  AND2X2 U56 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(n57) );
  AND2X2 U57 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(n58) );
  AND2X2 U58 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(n59) );
  AND2X2 U59 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(n60) );
  AND2X2 U60 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(n61) );
  AND2X2 U61 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(n62) );
  AND2X2 U62 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(n63) );
  AND2X2 U63 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n64) );
  AND2X2 U64 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(n65) );
  AND2X2 U65 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(n66) );
  XOR2X1 U68 ( .A(\SUMB[7][0] ), .B(n10), .Y(\A1[5] ) );
  XOR2X1 U69 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  XOR2X1 U70 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  XOR2X1 U71 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  XOR2X1 U72 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  XOR2X1 U73 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  XOR2X1 U74 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  XOR2X1 U75 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  XOR2X1 U76 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  XOR2X1 U77 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  XOR2X1 U78 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  XOR2X1 U79 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  XOR2X1 U80 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  XOR2X1 U81 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  XOR2X1 U82 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  XOR2X1 U83 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  XOR2X1 U84 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  XOR2X1 U85 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  XOR2X1 U86 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  XOR2X1 U87 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  XOR2X1 U88 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  XOR2X1 U89 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  XOR2X1 U90 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  XOR2X1 U91 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  XOR2X1 U92 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  XOR2X1 U93 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  XOR2X1 U94 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  XOR2X1 U95 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  XOR2X1 U96 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  XOR2X1 U97 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  XOR2X1 U98 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(\A1[36] ) );
  XOR2X1 U99 ( .A(\CARRYB[7][31] ), .B(TC), .Y(\A1[37] ) );
  XOR2X1 U100 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U101 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U102 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U103 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U104 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U105 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U106 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U107 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  XOR2X1 U108 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(\SUMB[1][8] ) );
  XOR2X1 U109 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Y(\SUMB[1][9] ) );
  XOR2X1 U110 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Y(\SUMB[1][10] ) );
  XOR2X1 U111 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U112 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Y(\SUMB[1][12] ) );
  XOR2X1 U113 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  XOR2X1 U114 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  XOR2X1 U115 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Y(\SUMB[1][15] ) );
  XOR2X1 U116 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Y(\SUMB[1][16] ) );
  XOR2X1 U117 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Y(\SUMB[1][17] ) );
  XOR2X1 U118 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Y(\SUMB[1][18] ) );
  XOR2X1 U119 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Y(\SUMB[1][19] ) );
  XOR2X1 U120 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Y(\SUMB[1][20] ) );
  XOR2X1 U121 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Y(\SUMB[1][21] ) );
  XOR2X1 U122 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Y(\SUMB[1][22] ) );
  XOR2X1 U123 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Y(\SUMB[1][23] ) );
  XOR2X1 U124 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Y(\SUMB[1][24] ) );
  XOR2X1 U125 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Y(\SUMB[1][25] ) );
  XOR2X1 U126 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Y(\SUMB[1][26] ) );
  XOR2X1 U127 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Y(\SUMB[1][27] ) );
  XOR2X1 U128 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Y(\SUMB[1][28] ) );
  XOR2X1 U129 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Y(\SUMB[1][29] ) );
  XOR2X1 U130 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Y(\SUMB[1][30] ) );
  MUX2X1 U171 ( .B(n129), .A(n130), .S(B[9]), .Y(\ab[7][9] ) );
  MUX2X1 U172 ( .B(n129), .A(n130), .S(B[8]), .Y(\ab[7][8] ) );
  MUX2X1 U173 ( .B(n129), .A(n130), .S(B[7]), .Y(\ab[7][7] ) );
  MUX2X1 U174 ( .B(n129), .A(n130), .S(B[6]), .Y(\ab[7][6] ) );
  MUX2X1 U175 ( .B(n129), .A(n130), .S(B[5]), .Y(\ab[7][5] ) );
  MUX2X1 U176 ( .B(n129), .A(n130), .S(B[4]), .Y(\ab[7][4] ) );
  MUX2X1 U177 ( .B(n129), .A(n130), .S(B[3]), .Y(\ab[7][3] ) );
  AND2X1 U178 ( .A(A[7]), .B(B[31]), .Y(\ab[7][31] ) );
  MUX2X1 U179 ( .B(n129), .A(n130), .S(B[30]), .Y(\ab[7][30] ) );
  MUX2X1 U180 ( .B(n129), .A(n130), .S(B[2]), .Y(\ab[7][2] ) );
  MUX2X1 U181 ( .B(n129), .A(n130), .S(B[29]), .Y(\ab[7][29] ) );
  MUX2X1 U182 ( .B(n129), .A(n130), .S(B[28]), .Y(\ab[7][28] ) );
  MUX2X1 U183 ( .B(n129), .A(n130), .S(B[27]), .Y(\ab[7][27] ) );
  MUX2X1 U184 ( .B(n129), .A(n130), .S(B[26]), .Y(\ab[7][26] ) );
  MUX2X1 U185 ( .B(n129), .A(n130), .S(B[25]), .Y(\ab[7][25] ) );
  MUX2X1 U186 ( .B(n129), .A(n130), .S(B[24]), .Y(\ab[7][24] ) );
  MUX2X1 U187 ( .B(n129), .A(n130), .S(B[23]), .Y(\ab[7][23] ) );
  MUX2X1 U188 ( .B(n129), .A(n130), .S(B[22]), .Y(\ab[7][22] ) );
  MUX2X1 U189 ( .B(n129), .A(n130), .S(B[21]), .Y(\ab[7][21] ) );
  MUX2X1 U190 ( .B(n129), .A(n130), .S(B[20]), .Y(\ab[7][20] ) );
  MUX2X1 U191 ( .B(n129), .A(n130), .S(B[1]), .Y(\ab[7][1] ) );
  MUX2X1 U192 ( .B(n129), .A(n130), .S(B[19]), .Y(\ab[7][19] ) );
  MUX2X1 U193 ( .B(n129), .A(n130), .S(B[18]), .Y(\ab[7][18] ) );
  MUX2X1 U194 ( .B(n129), .A(n130), .S(B[17]), .Y(\ab[7][17] ) );
  MUX2X1 U195 ( .B(n129), .A(n130), .S(B[16]), .Y(\ab[7][16] ) );
  MUX2X1 U196 ( .B(n129), .A(n130), .S(B[15]), .Y(\ab[7][15] ) );
  MUX2X1 U197 ( .B(n129), .A(n130), .S(B[14]), .Y(\ab[7][14] ) );
  MUX2X1 U198 ( .B(n129), .A(n130), .S(B[13]), .Y(\ab[7][13] ) );
  MUX2X1 U199 ( .B(n129), .A(n130), .S(B[12]), .Y(\ab[7][12] ) );
  MUX2X1 U200 ( .B(n129), .A(n130), .S(B[11]), .Y(\ab[7][11] ) );
  MUX2X1 U201 ( .B(n129), .A(n130), .S(B[10]), .Y(\ab[7][10] ) );
  MUX2X1 U202 ( .B(n129), .A(n130), .S(B[0]), .Y(\ab[7][0] ) );
  NOR2X1 U203 ( .A(n154), .B(n128), .Y(\ab[6][9] ) );
  NOR2X1 U204 ( .A(n153), .B(n128), .Y(\ab[6][8] ) );
  NOR2X1 U205 ( .A(n114), .B(n128), .Y(\ab[6][7] ) );
  NOR2X1 U206 ( .A(n115), .B(n128), .Y(\ab[6][6] ) );
  NOR2X1 U207 ( .A(n116), .B(n128), .Y(\ab[6][5] ) );
  NOR2X1 U208 ( .A(n117), .B(n128), .Y(\ab[6][4] ) );
  NOR2X1 U209 ( .A(n118), .B(n128), .Y(\ab[6][3] ) );
  MUX2X1 U210 ( .B(n110), .A(n111), .S(A[6]), .Y(\ab[6][31] ) );
  NOR2X1 U211 ( .A(n151), .B(n128), .Y(\ab[6][30] ) );
  NOR2X1 U212 ( .A(n119), .B(n128), .Y(\ab[6][2] ) );
  NOR2X1 U213 ( .A(n150), .B(n128), .Y(\ab[6][29] ) );
  NOR2X1 U214 ( .A(n149), .B(n128), .Y(\ab[6][28] ) );
  NOR2X1 U215 ( .A(n148), .B(n128), .Y(\ab[6][27] ) );
  NOR2X1 U216 ( .A(n147), .B(n128), .Y(\ab[6][26] ) );
  NOR2X1 U217 ( .A(n146), .B(n128), .Y(\ab[6][25] ) );
  NOR2X1 U218 ( .A(n145), .B(n128), .Y(\ab[6][24] ) );
  NOR2X1 U219 ( .A(n144), .B(n128), .Y(\ab[6][23] ) );
  NOR2X1 U220 ( .A(n143), .B(n128), .Y(\ab[6][22] ) );
  NOR2X1 U221 ( .A(n142), .B(n128), .Y(\ab[6][21] ) );
  NOR2X1 U222 ( .A(n141), .B(n128), .Y(\ab[6][20] ) );
  NOR2X1 U223 ( .A(n120), .B(n128), .Y(\ab[6][1] ) );
  NOR2X1 U224 ( .A(n140), .B(n128), .Y(\ab[6][19] ) );
  NOR2X1 U225 ( .A(n139), .B(n128), .Y(\ab[6][18] ) );
  NOR2X1 U226 ( .A(n138), .B(n128), .Y(\ab[6][17] ) );
  NOR2X1 U227 ( .A(n137), .B(n128), .Y(\ab[6][16] ) );
  NOR2X1 U228 ( .A(n136), .B(n128), .Y(\ab[6][15] ) );
  NOR2X1 U229 ( .A(n135), .B(n128), .Y(\ab[6][14] ) );
  NOR2X1 U230 ( .A(n134), .B(n128), .Y(\ab[6][13] ) );
  NOR2X1 U231 ( .A(n133), .B(n128), .Y(\ab[6][12] ) );
  NOR2X1 U232 ( .A(n132), .B(n128), .Y(\ab[6][11] ) );
  NOR2X1 U233 ( .A(n131), .B(n128), .Y(\ab[6][10] ) );
  NOR2X1 U234 ( .A(n122), .B(n128), .Y(\ab[6][0] ) );
  NOR2X1 U235 ( .A(n154), .B(n127), .Y(\ab[5][9] ) );
  NOR2X1 U236 ( .A(n153), .B(n127), .Y(\ab[5][8] ) );
  NOR2X1 U237 ( .A(n114), .B(n127), .Y(\ab[5][7] ) );
  NOR2X1 U238 ( .A(n115), .B(n127), .Y(\ab[5][6] ) );
  NOR2X1 U239 ( .A(n116), .B(n127), .Y(\ab[5][5] ) );
  NOR2X1 U240 ( .A(n117), .B(n127), .Y(\ab[5][4] ) );
  NOR2X1 U241 ( .A(n118), .B(n127), .Y(\ab[5][3] ) );
  MUX2X1 U242 ( .B(n110), .A(n111), .S(A[5]), .Y(\ab[5][31] ) );
  NOR2X1 U243 ( .A(n151), .B(n127), .Y(\ab[5][30] ) );
  NOR2X1 U244 ( .A(n119), .B(n127), .Y(\ab[5][2] ) );
  NOR2X1 U245 ( .A(n150), .B(n127), .Y(\ab[5][29] ) );
  NOR2X1 U246 ( .A(n149), .B(n127), .Y(\ab[5][28] ) );
  NOR2X1 U247 ( .A(n148), .B(n127), .Y(\ab[5][27] ) );
  NOR2X1 U248 ( .A(n147), .B(n127), .Y(\ab[5][26] ) );
  NOR2X1 U249 ( .A(n146), .B(n127), .Y(\ab[5][25] ) );
  NOR2X1 U250 ( .A(n145), .B(n127), .Y(\ab[5][24] ) );
  NOR2X1 U251 ( .A(n144), .B(n127), .Y(\ab[5][23] ) );
  NOR2X1 U252 ( .A(n143), .B(n127), .Y(\ab[5][22] ) );
  NOR2X1 U253 ( .A(n142), .B(n127), .Y(\ab[5][21] ) );
  NOR2X1 U254 ( .A(n141), .B(n127), .Y(\ab[5][20] ) );
  NOR2X1 U255 ( .A(n120), .B(n127), .Y(\ab[5][1] ) );
  NOR2X1 U256 ( .A(n140), .B(n127), .Y(\ab[5][19] ) );
  NOR2X1 U257 ( .A(n139), .B(n127), .Y(\ab[5][18] ) );
  NOR2X1 U258 ( .A(n138), .B(n127), .Y(\ab[5][17] ) );
  NOR2X1 U259 ( .A(n137), .B(n127), .Y(\ab[5][16] ) );
  NOR2X1 U260 ( .A(n136), .B(n127), .Y(\ab[5][15] ) );
  NOR2X1 U261 ( .A(n135), .B(n127), .Y(\ab[5][14] ) );
  NOR2X1 U262 ( .A(n134), .B(n127), .Y(\ab[5][13] ) );
  NOR2X1 U263 ( .A(n133), .B(n127), .Y(\ab[5][12] ) );
  NOR2X1 U264 ( .A(n132), .B(n127), .Y(\ab[5][11] ) );
  NOR2X1 U265 ( .A(n131), .B(n127), .Y(\ab[5][10] ) );
  NOR2X1 U266 ( .A(n122), .B(n127), .Y(\ab[5][0] ) );
  NOR2X1 U267 ( .A(n154), .B(n126), .Y(\ab[4][9] ) );
  NOR2X1 U268 ( .A(n153), .B(n126), .Y(\ab[4][8] ) );
  NOR2X1 U269 ( .A(n114), .B(n126), .Y(\ab[4][7] ) );
  NOR2X1 U270 ( .A(n115), .B(n126), .Y(\ab[4][6] ) );
  NOR2X1 U271 ( .A(n116), .B(n126), .Y(\ab[4][5] ) );
  NOR2X1 U272 ( .A(n117), .B(n126), .Y(\ab[4][4] ) );
  NOR2X1 U273 ( .A(n118), .B(n126), .Y(\ab[4][3] ) );
  MUX2X1 U274 ( .B(n110), .A(n111), .S(A[4]), .Y(\ab[4][31] ) );
  NOR2X1 U275 ( .A(n151), .B(n126), .Y(\ab[4][30] ) );
  NOR2X1 U276 ( .A(n119), .B(n126), .Y(\ab[4][2] ) );
  NOR2X1 U277 ( .A(n150), .B(n126), .Y(\ab[4][29] ) );
  NOR2X1 U278 ( .A(n149), .B(n126), .Y(\ab[4][28] ) );
  NOR2X1 U279 ( .A(n148), .B(n126), .Y(\ab[4][27] ) );
  NOR2X1 U280 ( .A(n147), .B(n126), .Y(\ab[4][26] ) );
  NOR2X1 U281 ( .A(n146), .B(n126), .Y(\ab[4][25] ) );
  NOR2X1 U282 ( .A(n145), .B(n126), .Y(\ab[4][24] ) );
  NOR2X1 U283 ( .A(n144), .B(n126), .Y(\ab[4][23] ) );
  NOR2X1 U284 ( .A(n143), .B(n126), .Y(\ab[4][22] ) );
  NOR2X1 U285 ( .A(n142), .B(n126), .Y(\ab[4][21] ) );
  NOR2X1 U286 ( .A(n141), .B(n126), .Y(\ab[4][20] ) );
  NOR2X1 U287 ( .A(n120), .B(n126), .Y(\ab[4][1] ) );
  NOR2X1 U288 ( .A(n140), .B(n126), .Y(\ab[4][19] ) );
  NOR2X1 U289 ( .A(n139), .B(n126), .Y(\ab[4][18] ) );
  NOR2X1 U290 ( .A(n138), .B(n126), .Y(\ab[4][17] ) );
  NOR2X1 U291 ( .A(n137), .B(n126), .Y(\ab[4][16] ) );
  NOR2X1 U292 ( .A(n136), .B(n126), .Y(\ab[4][15] ) );
  NOR2X1 U293 ( .A(n135), .B(n126), .Y(\ab[4][14] ) );
  NOR2X1 U294 ( .A(n134), .B(n126), .Y(\ab[4][13] ) );
  NOR2X1 U295 ( .A(n133), .B(n126), .Y(\ab[4][12] ) );
  NOR2X1 U296 ( .A(n132), .B(n126), .Y(\ab[4][11] ) );
  NOR2X1 U297 ( .A(n131), .B(n126), .Y(\ab[4][10] ) );
  NOR2X1 U298 ( .A(n122), .B(n126), .Y(\ab[4][0] ) );
  NOR2X1 U299 ( .A(n154), .B(n125), .Y(\ab[3][9] ) );
  NOR2X1 U300 ( .A(n153), .B(n125), .Y(\ab[3][8] ) );
  NOR2X1 U301 ( .A(n114), .B(n125), .Y(\ab[3][7] ) );
  NOR2X1 U302 ( .A(n115), .B(n125), .Y(\ab[3][6] ) );
  NOR2X1 U303 ( .A(n116), .B(n125), .Y(\ab[3][5] ) );
  NOR2X1 U304 ( .A(n117), .B(n125), .Y(\ab[3][4] ) );
  NOR2X1 U305 ( .A(n118), .B(n125), .Y(\ab[3][3] ) );
  MUX2X1 U306 ( .B(n110), .A(n111), .S(A[3]), .Y(\ab[3][31] ) );
  NOR2X1 U307 ( .A(n151), .B(n125), .Y(\ab[3][30] ) );
  NOR2X1 U308 ( .A(n119), .B(n125), .Y(\ab[3][2] ) );
  NOR2X1 U309 ( .A(n150), .B(n125), .Y(\ab[3][29] ) );
  NOR2X1 U310 ( .A(n149), .B(n125), .Y(\ab[3][28] ) );
  NOR2X1 U311 ( .A(n148), .B(n125), .Y(\ab[3][27] ) );
  NOR2X1 U312 ( .A(n147), .B(n125), .Y(\ab[3][26] ) );
  NOR2X1 U313 ( .A(n146), .B(n125), .Y(\ab[3][25] ) );
  NOR2X1 U314 ( .A(n145), .B(n125), .Y(\ab[3][24] ) );
  NOR2X1 U315 ( .A(n144), .B(n125), .Y(\ab[3][23] ) );
  NOR2X1 U316 ( .A(n143), .B(n125), .Y(\ab[3][22] ) );
  NOR2X1 U317 ( .A(n142), .B(n125), .Y(\ab[3][21] ) );
  NOR2X1 U318 ( .A(n141), .B(n125), .Y(\ab[3][20] ) );
  NOR2X1 U319 ( .A(n120), .B(n125), .Y(\ab[3][1] ) );
  NOR2X1 U320 ( .A(n140), .B(n125), .Y(\ab[3][19] ) );
  NOR2X1 U321 ( .A(n139), .B(n125), .Y(\ab[3][18] ) );
  NOR2X1 U322 ( .A(n138), .B(n125), .Y(\ab[3][17] ) );
  NOR2X1 U323 ( .A(n137), .B(n125), .Y(\ab[3][16] ) );
  NOR2X1 U324 ( .A(n136), .B(n125), .Y(\ab[3][15] ) );
  NOR2X1 U325 ( .A(n135), .B(n125), .Y(\ab[3][14] ) );
  NOR2X1 U326 ( .A(n134), .B(n125), .Y(\ab[3][13] ) );
  NOR2X1 U327 ( .A(n133), .B(n125), .Y(\ab[3][12] ) );
  NOR2X1 U328 ( .A(n132), .B(n125), .Y(\ab[3][11] ) );
  NOR2X1 U329 ( .A(n131), .B(n125), .Y(\ab[3][10] ) );
  NOR2X1 U330 ( .A(n122), .B(n125), .Y(\ab[3][0] ) );
  NOR2X1 U331 ( .A(n154), .B(n121), .Y(\ab[2][9] ) );
  NOR2X1 U332 ( .A(n153), .B(n121), .Y(\ab[2][8] ) );
  NOR2X1 U333 ( .A(n114), .B(n121), .Y(\ab[2][7] ) );
  NOR2X1 U334 ( .A(n115), .B(n121), .Y(\ab[2][6] ) );
  NOR2X1 U335 ( .A(n116), .B(n121), .Y(\ab[2][5] ) );
  NOR2X1 U336 ( .A(n117), .B(n121), .Y(\ab[2][4] ) );
  NOR2X1 U337 ( .A(n118), .B(n121), .Y(\ab[2][3] ) );
  MUX2X1 U338 ( .B(n110), .A(n111), .S(A[2]), .Y(\ab[2][31] ) );
  NOR2X1 U339 ( .A(n151), .B(n121), .Y(\ab[2][30] ) );
  NOR2X1 U340 ( .A(n119), .B(n121), .Y(\ab[2][2] ) );
  NOR2X1 U341 ( .A(n150), .B(n121), .Y(\ab[2][29] ) );
  NOR2X1 U342 ( .A(n149), .B(n121), .Y(\ab[2][28] ) );
  NOR2X1 U343 ( .A(n148), .B(n121), .Y(\ab[2][27] ) );
  NOR2X1 U344 ( .A(n147), .B(n121), .Y(\ab[2][26] ) );
  NOR2X1 U345 ( .A(n146), .B(n121), .Y(\ab[2][25] ) );
  NOR2X1 U346 ( .A(n145), .B(n121), .Y(\ab[2][24] ) );
  NOR2X1 U347 ( .A(n144), .B(n121), .Y(\ab[2][23] ) );
  NOR2X1 U348 ( .A(n143), .B(n121), .Y(\ab[2][22] ) );
  NOR2X1 U349 ( .A(n142), .B(n121), .Y(\ab[2][21] ) );
  NOR2X1 U350 ( .A(n141), .B(n121), .Y(\ab[2][20] ) );
  NOR2X1 U351 ( .A(n120), .B(n121), .Y(\ab[2][1] ) );
  NOR2X1 U352 ( .A(n140), .B(n121), .Y(\ab[2][19] ) );
  NOR2X1 U353 ( .A(n139), .B(n121), .Y(\ab[2][18] ) );
  NOR2X1 U354 ( .A(n138), .B(n121), .Y(\ab[2][17] ) );
  NOR2X1 U355 ( .A(n137), .B(n121), .Y(\ab[2][16] ) );
  NOR2X1 U356 ( .A(n136), .B(n121), .Y(\ab[2][15] ) );
  NOR2X1 U357 ( .A(n135), .B(n121), .Y(\ab[2][14] ) );
  NOR2X1 U358 ( .A(n134), .B(n121), .Y(\ab[2][13] ) );
  NOR2X1 U359 ( .A(n133), .B(n121), .Y(\ab[2][12] ) );
  NOR2X1 U360 ( .A(n132), .B(n121), .Y(\ab[2][11] ) );
  NOR2X1 U361 ( .A(n131), .B(n121), .Y(\ab[2][10] ) );
  NOR2X1 U362 ( .A(n122), .B(n121), .Y(\ab[2][0] ) );
  NOR2X1 U363 ( .A(n154), .B(n124), .Y(\ab[1][9] ) );
  NOR2X1 U364 ( .A(n153), .B(n124), .Y(\ab[1][8] ) );
  NOR2X1 U365 ( .A(n114), .B(n124), .Y(\ab[1][7] ) );
  NOR2X1 U366 ( .A(n115), .B(n124), .Y(\ab[1][6] ) );
  NOR2X1 U367 ( .A(n116), .B(n124), .Y(\ab[1][5] ) );
  NOR2X1 U368 ( .A(n117), .B(n124), .Y(\ab[1][4] ) );
  NOR2X1 U369 ( .A(n118), .B(n124), .Y(\ab[1][3] ) );
  MUX2X1 U370 ( .B(n110), .A(n111), .S(A[1]), .Y(\ab[1][31] ) );
  NOR2X1 U371 ( .A(n151), .B(n124), .Y(\ab[1][30] ) );
  NOR2X1 U372 ( .A(n119), .B(n124), .Y(\ab[1][2] ) );
  NOR2X1 U373 ( .A(n150), .B(n124), .Y(\ab[1][29] ) );
  NOR2X1 U374 ( .A(n149), .B(n124), .Y(\ab[1][28] ) );
  NOR2X1 U375 ( .A(n148), .B(n124), .Y(\ab[1][27] ) );
  NOR2X1 U376 ( .A(n147), .B(n124), .Y(\ab[1][26] ) );
  NOR2X1 U377 ( .A(n146), .B(n124), .Y(\ab[1][25] ) );
  NOR2X1 U378 ( .A(n145), .B(n124), .Y(\ab[1][24] ) );
  NOR2X1 U379 ( .A(n144), .B(n124), .Y(\ab[1][23] ) );
  NOR2X1 U380 ( .A(n143), .B(n124), .Y(\ab[1][22] ) );
  NOR2X1 U381 ( .A(n142), .B(n124), .Y(\ab[1][21] ) );
  NOR2X1 U382 ( .A(n141), .B(n124), .Y(\ab[1][20] ) );
  NOR2X1 U383 ( .A(n120), .B(n124), .Y(\ab[1][1] ) );
  NOR2X1 U384 ( .A(n140), .B(n124), .Y(\ab[1][19] ) );
  NOR2X1 U385 ( .A(n139), .B(n124), .Y(\ab[1][18] ) );
  NOR2X1 U386 ( .A(n138), .B(n124), .Y(\ab[1][17] ) );
  NOR2X1 U387 ( .A(n137), .B(n124), .Y(\ab[1][16] ) );
  NOR2X1 U388 ( .A(n136), .B(n124), .Y(\ab[1][15] ) );
  NOR2X1 U389 ( .A(n135), .B(n124), .Y(\ab[1][14] ) );
  NOR2X1 U390 ( .A(n134), .B(n124), .Y(\ab[1][13] ) );
  NOR2X1 U391 ( .A(n133), .B(n124), .Y(\ab[1][12] ) );
  NOR2X1 U392 ( .A(n132), .B(n124), .Y(\ab[1][11] ) );
  NOR2X1 U393 ( .A(n131), .B(n124), .Y(\ab[1][10] ) );
  NOR2X1 U394 ( .A(n122), .B(n124), .Y(\ab[1][0] ) );
  NOR2X1 U395 ( .A(n154), .B(n123), .Y(\ab[0][9] ) );
  NOR2X1 U396 ( .A(n153), .B(n123), .Y(\ab[0][8] ) );
  NOR2X1 U397 ( .A(n114), .B(n123), .Y(\ab[0][7] ) );
  NOR2X1 U398 ( .A(n115), .B(n123), .Y(\ab[0][6] ) );
  NOR2X1 U399 ( .A(n116), .B(n123), .Y(\ab[0][5] ) );
  NOR2X1 U400 ( .A(n117), .B(n123), .Y(\ab[0][4] ) );
  NOR2X1 U401 ( .A(n118), .B(n123), .Y(\ab[0][3] ) );
  MUX2X1 U402 ( .B(n110), .A(n111), .S(A[0]), .Y(\ab[0][31] ) );
  NAND2X1 U403 ( .A(B[31]), .B(n155), .Y(n111) );
  NOR2X1 U404 ( .A(n151), .B(n123), .Y(\ab[0][30] ) );
  NOR2X1 U405 ( .A(n119), .B(n123), .Y(\ab[0][2] ) );
  NOR2X1 U406 ( .A(n150), .B(n123), .Y(\ab[0][29] ) );
  NOR2X1 U407 ( .A(n149), .B(n123), .Y(\ab[0][28] ) );
  NOR2X1 U408 ( .A(n148), .B(n123), .Y(\ab[0][27] ) );
  NOR2X1 U409 ( .A(n147), .B(n123), .Y(\ab[0][26] ) );
  NOR2X1 U410 ( .A(n146), .B(n123), .Y(\ab[0][25] ) );
  NOR2X1 U411 ( .A(n145), .B(n123), .Y(\ab[0][24] ) );
  NOR2X1 U412 ( .A(n144), .B(n123), .Y(\ab[0][23] ) );
  NOR2X1 U413 ( .A(n143), .B(n123), .Y(\ab[0][22] ) );
  NOR2X1 U414 ( .A(n142), .B(n123), .Y(\ab[0][21] ) );
  NOR2X1 U415 ( .A(n141), .B(n123), .Y(\ab[0][20] ) );
  NOR2X1 U416 ( .A(n120), .B(n123), .Y(\ab[0][1] ) );
  NOR2X1 U417 ( .A(n140), .B(n123), .Y(\ab[0][19] ) );
  NOR2X1 U418 ( .A(n139), .B(n123), .Y(\ab[0][18] ) );
  NOR2X1 U419 ( .A(n138), .B(n123), .Y(\ab[0][17] ) );
  NOR2X1 U420 ( .A(n137), .B(n123), .Y(\ab[0][16] ) );
  NOR2X1 U421 ( .A(n136), .B(n123), .Y(\ab[0][15] ) );
  NOR2X1 U422 ( .A(n135), .B(n123), .Y(\ab[0][14] ) );
  NOR2X1 U423 ( .A(n134), .B(n123), .Y(\ab[0][13] ) );
  NOR2X1 U424 ( .A(n133), .B(n123), .Y(\ab[0][12] ) );
  NOR2X1 U425 ( .A(n132), .B(n123), .Y(\ab[0][11] ) );
  NOR2X1 U426 ( .A(n131), .B(n123), .Y(\ab[0][10] ) );
  NAND2X1 U427 ( .A(B[31]), .B(TC), .Y(n110) );
  NOR2X1 U428 ( .A(B[31]), .B(n155), .Y(QB) );
  NOR2X1 U429 ( .A(A[7]), .B(n155), .Y(QA) );
  NOR2X1 U430 ( .A(n122), .B(n123), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_41 FS_1 ( .A({\A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n9, n8, n7, 
        n6, n5, n4, n3, \A2[30] , n45, n54, n46, n55, n47, n56, n48, n57, n49, 
        n58, n50, n59, n51, n60, n52, n61, n53, n62, n63, n66, n64, n65, n43, 
        n44, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  INVX2 U131 ( .A(B[7]), .Y(n114) );
  INVX2 U132 ( .A(B[6]), .Y(n115) );
  INVX2 U133 ( .A(B[5]), .Y(n116) );
  INVX2 U134 ( .A(B[4]), .Y(n117) );
  INVX2 U135 ( .A(B[3]), .Y(n118) );
  INVX2 U136 ( .A(B[2]), .Y(n119) );
  INVX2 U137 ( .A(B[1]), .Y(n120) );
  INVX2 U138 ( .A(A[2]), .Y(n121) );
  INVX2 U139 ( .A(B[0]), .Y(n122) );
  INVX2 U140 ( .A(A[0]), .Y(n123) );
  INVX2 U141 ( .A(A[1]), .Y(n124) );
  INVX2 U142 ( .A(A[3]), .Y(n125) );
  INVX2 U143 ( .A(A[4]), .Y(n126) );
  INVX2 U144 ( .A(A[5]), .Y(n127) );
  INVX2 U145 ( .A(A[6]), .Y(n128) );
  INVX2 U146 ( .A(n10), .Y(n129) );
  INVX2 U147 ( .A(n11), .Y(n130) );
  INVX2 U148 ( .A(B[10]), .Y(n131) );
  INVX2 U149 ( .A(B[11]), .Y(n132) );
  INVX2 U150 ( .A(B[12]), .Y(n133) );
  INVX2 U151 ( .A(B[13]), .Y(n134) );
  INVX2 U152 ( .A(B[14]), .Y(n135) );
  INVX2 U153 ( .A(B[15]), .Y(n136) );
  INVX2 U154 ( .A(B[16]), .Y(n137) );
  INVX2 U155 ( .A(B[17]), .Y(n138) );
  INVX2 U156 ( .A(B[18]), .Y(n139) );
  INVX2 U157 ( .A(B[19]), .Y(n140) );
  INVX2 U158 ( .A(B[20]), .Y(n141) );
  INVX2 U159 ( .A(B[21]), .Y(n142) );
  INVX2 U160 ( .A(B[22]), .Y(n143) );
  INVX2 U161 ( .A(B[23]), .Y(n144) );
  INVX2 U162 ( .A(B[24]), .Y(n145) );
  INVX2 U163 ( .A(B[25]), .Y(n146) );
  INVX2 U164 ( .A(B[26]), .Y(n147) );
  INVX2 U165 ( .A(B[27]), .Y(n148) );
  INVX2 U166 ( .A(B[28]), .Y(n149) );
  INVX2 U167 ( .A(B[29]), .Y(n150) );
  INVX2 U168 ( .A(B[30]), .Y(n151) );
  INVX2 U169 ( .A(n110), .Y(n152) );
  INVX2 U170 ( .A(B[8]), .Y(n153) );
  INVX2 U431 ( .A(B[9]), .Y(n154) );
  INVX2 U432 ( .A(TC), .Y(n155) );
endmodule


module CannyEdge_DW01_cmp2_4 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188;

  MUX2X1 U63 ( .B(n63), .A(n64), .S(B[31]), .Y(GE_GT) );
  MUX2X1 U64 ( .B(TC), .A(n65), .S(A[31]), .Y(n64) );
  NOR2X1 U65 ( .A(n66), .B(n167), .Y(n65) );
  MUX2X1 U66 ( .B(n67), .A(n188), .S(A[31]), .Y(n63) );
  NAND2X1 U67 ( .A(n66), .B(n167), .Y(n67) );
  OAI21X1 U68 ( .A(A[29]), .B(n147), .C(n68), .Y(n66) );
  OAI21X1 U69 ( .A(B[29]), .B(n168), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(A[28]), .B(n146), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(B[28]), .B(n169), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(A[27]), .B(n145), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(B[27]), .B(n170), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(A[26]), .B(n144), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(B[26]), .B(n171), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(A[25]), .B(n143), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(B[25]), .B(n172), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(A[24]), .B(n142), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(B[24]), .B(n173), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(A[23]), .B(n141), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(B[23]), .B(n174), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(A[22]), .B(n140), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(B[22]), .B(n175), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(A[21]), .B(n139), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(B[21]), .B(n176), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(A[20]), .B(n138), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(B[20]), .B(n177), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(A[19]), .B(n137), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(B[19]), .B(n178), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(A[18]), .B(n136), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(B[18]), .B(n179), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(A[17]), .B(n135), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(B[17]), .B(n180), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(A[16]), .B(n148), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(B[16]), .B(n181), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(A[15]), .B(n149), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(B[15]), .B(n182), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(A[14]), .B(n150), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(B[14]), .B(n183), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(A[13]), .B(n151), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(B[13]), .B(n184), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(A[12]), .B(n152), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(B[12]), .B(n185), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(A[11]), .B(n153), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(B[11]), .B(n186), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(A[10]), .B(n154), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(B[10]), .B(n187), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(A[9]), .B(n155), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(B[9]), .B(n165), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(A[8]), .B(n156), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(B[8]), .B(n166), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(A[7]), .B(n157), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(B[7]), .B(n134), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(A[6]), .B(n158), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(B[6]), .B(n133), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(A[5]), .B(n159), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(B[5]), .B(n132), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(A[4]), .B(n160), .C(n118), .Y(n117) );
  AOI21X1 U119 ( .A(B[4]), .B(n131), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(A[3]), .B(n161), .C(n120), .Y(n119) );
  OAI21X1 U121 ( .A(B[3]), .B(n130), .C(n121), .Y(n120) );
  AOI21X1 U122 ( .A(A[2]), .B(n162), .C(n122), .Y(n121) );
  AOI21X1 U123 ( .A(B[2]), .B(n129), .C(n123), .Y(n122) );
  OAI21X1 U124 ( .A(A[1]), .B(n163), .C(n124), .Y(n123) );
  OAI21X1 U125 ( .A(B[1]), .B(n128), .C(n125), .Y(n124) );
  AOI21X1 U126 ( .A(A[0]), .B(n164), .C(n126), .Y(n125) );
  AOI21X1 U127 ( .A(B[0]), .B(n127), .C(LEQ), .Y(n126) );
  INVX2 U1 ( .A(A[0]), .Y(n127) );
  INVX2 U2 ( .A(A[1]), .Y(n128) );
  INVX2 U3 ( .A(A[2]), .Y(n129) );
  INVX2 U4 ( .A(A[3]), .Y(n130) );
  INVX2 U5 ( .A(A[4]), .Y(n131) );
  INVX2 U6 ( .A(A[5]), .Y(n132) );
  INVX2 U7 ( .A(A[6]), .Y(n133) );
  INVX2 U8 ( .A(A[7]), .Y(n134) );
  INVX2 U9 ( .A(B[17]), .Y(n135) );
  INVX2 U10 ( .A(B[18]), .Y(n136) );
  INVX2 U11 ( .A(B[19]), .Y(n137) );
  INVX2 U12 ( .A(B[20]), .Y(n138) );
  INVX2 U13 ( .A(B[21]), .Y(n139) );
  INVX2 U14 ( .A(B[22]), .Y(n140) );
  INVX2 U15 ( .A(B[23]), .Y(n141) );
  INVX2 U16 ( .A(B[24]), .Y(n142) );
  INVX2 U17 ( .A(B[25]), .Y(n143) );
  INVX2 U18 ( .A(B[26]), .Y(n144) );
  INVX2 U19 ( .A(B[27]), .Y(n145) );
  INVX2 U20 ( .A(B[28]), .Y(n146) );
  INVX2 U21 ( .A(B[29]), .Y(n147) );
  INVX2 U22 ( .A(B[16]), .Y(n148) );
  INVX2 U23 ( .A(B[15]), .Y(n149) );
  INVX2 U24 ( .A(B[14]), .Y(n150) );
  INVX2 U25 ( .A(B[13]), .Y(n151) );
  INVX2 U26 ( .A(B[12]), .Y(n152) );
  INVX2 U27 ( .A(B[11]), .Y(n153) );
  INVX2 U28 ( .A(B[10]), .Y(n154) );
  INVX2 U29 ( .A(B[9]), .Y(n155) );
  INVX2 U30 ( .A(B[8]), .Y(n156) );
  INVX2 U31 ( .A(B[7]), .Y(n157) );
  INVX2 U32 ( .A(B[6]), .Y(n158) );
  INVX2 U33 ( .A(B[5]), .Y(n159) );
  INVX2 U34 ( .A(B[4]), .Y(n160) );
  INVX2 U35 ( .A(B[3]), .Y(n161) );
  INVX2 U36 ( .A(B[2]), .Y(n162) );
  INVX2 U37 ( .A(B[1]), .Y(n163) );
  INVX2 U38 ( .A(B[0]), .Y(n164) );
  INVX2 U39 ( .A(A[9]), .Y(n165) );
  INVX2 U40 ( .A(A[8]), .Y(n166) );
  INVX2 U41 ( .A(A[30]), .Y(n167) );
  INVX2 U42 ( .A(A[29]), .Y(n168) );
  INVX2 U43 ( .A(A[28]), .Y(n169) );
  INVX2 U44 ( .A(A[27]), .Y(n170) );
  INVX2 U45 ( .A(A[26]), .Y(n171) );
  INVX2 U46 ( .A(A[25]), .Y(n172) );
  INVX2 U47 ( .A(A[24]), .Y(n173) );
  INVX2 U48 ( .A(A[23]), .Y(n174) );
  INVX2 U49 ( .A(A[22]), .Y(n175) );
  INVX2 U50 ( .A(A[21]), .Y(n176) );
  INVX2 U51 ( .A(A[20]), .Y(n177) );
  INVX2 U52 ( .A(A[19]), .Y(n178) );
  INVX2 U53 ( .A(A[18]), .Y(n179) );
  INVX2 U54 ( .A(A[17]), .Y(n180) );
  INVX2 U55 ( .A(A[16]), .Y(n181) );
  INVX2 U56 ( .A(A[15]), .Y(n182) );
  INVX2 U57 ( .A(A[14]), .Y(n183) );
  INVX2 U58 ( .A(A[13]), .Y(n184) );
  INVX2 U59 ( .A(A[12]), .Y(n185) );
  INVX2 U60 ( .A(A[11]), .Y(n186) );
  INVX2 U61 ( .A(A[10]), .Y(n187) );
  INVX2 U62 ( .A(TC), .Y(n188) );
endmodule


module CannyEdge_DW01_add_42 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n141, n142, n143, n144, n145, n146, n147,
         n148, n149;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U31 ( .A(n30), .B(n31), .Y(SUM[9]) );
  NOR2X1 U32 ( .A(n130), .B(n32), .Y(n31) );
  XOR2X1 U33 ( .A(n34), .B(n134), .Y(SUM[8]) );
  NAND2X1 U34 ( .A(n133), .B(n35), .Y(n34) );
  XOR2X1 U35 ( .A(n37), .B(n38), .Y(SUM[7]) );
  XOR2X1 U36 ( .A(n135), .B(B[7]), .Y(n38) );
  OAI21X1 U37 ( .A(B[6]), .B(A[6]), .C(n37), .Y(n39) );
  XOR2X1 U38 ( .A(n40), .B(n41), .Y(SUM[29]) );
  XOR2X1 U39 ( .A(B[29]), .B(A[29]), .Y(n41) );
  OAI21X1 U40 ( .A(n42), .B(n43), .C(n44), .Y(n40) );
  XOR2X1 U41 ( .A(n45), .B(n43), .Y(SUM[28]) );
  AOI21X1 U42 ( .A(n137), .B(n46), .C(n47), .Y(n43) );
  NAND2X1 U43 ( .A(n136), .B(n44), .Y(n45) );
  NAND2X1 U44 ( .A(B[28]), .B(A[28]), .Y(n44) );
  NOR2X1 U45 ( .A(B[28]), .B(A[28]), .Y(n42) );
  XOR2X1 U46 ( .A(n46), .B(n49), .Y(SUM[27]) );
  NOR2X1 U47 ( .A(n47), .B(n48), .Y(n49) );
  NOR2X1 U48 ( .A(B[27]), .B(A[27]), .Y(n48) );
  AND2X1 U49 ( .A(B[27]), .B(A[27]), .Y(n47) );
  OAI21X1 U50 ( .A(n50), .B(n51), .C(n52), .Y(n46) );
  XOR2X1 U51 ( .A(n53), .B(n51), .Y(SUM[26]) );
  AOI21X1 U52 ( .A(n139), .B(n54), .C(n55), .Y(n51) );
  NAND2X1 U53 ( .A(n138), .B(n52), .Y(n53) );
  NAND2X1 U54 ( .A(B[26]), .B(A[26]), .Y(n52) );
  NOR2X1 U55 ( .A(B[26]), .B(A[26]), .Y(n50) );
  XOR2X1 U56 ( .A(n54), .B(n57), .Y(SUM[25]) );
  NOR2X1 U57 ( .A(n55), .B(n56), .Y(n57) );
  NOR2X1 U58 ( .A(B[25]), .B(A[25]), .Y(n56) );
  AND2X1 U59 ( .A(B[25]), .B(A[25]), .Y(n55) );
  OAI21X1 U60 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  XOR2X1 U61 ( .A(n61), .B(n59), .Y(SUM[24]) );
  AOI21X1 U62 ( .A(n143), .B(n62), .C(n63), .Y(n59) );
  NAND2X1 U63 ( .A(n142), .B(n60), .Y(n61) );
  NAND2X1 U64 ( .A(B[24]), .B(A[24]), .Y(n60) );
  NOR2X1 U65 ( .A(B[24]), .B(A[24]), .Y(n58) );
  XOR2X1 U66 ( .A(n62), .B(n65), .Y(SUM[23]) );
  NOR2X1 U67 ( .A(n63), .B(n64), .Y(n65) );
  NOR2X1 U68 ( .A(B[23]), .B(A[23]), .Y(n64) );
  AND2X1 U69 ( .A(B[23]), .B(A[23]), .Y(n63) );
  OAI21X1 U70 ( .A(n66), .B(n67), .C(n68), .Y(n62) );
  XOR2X1 U71 ( .A(n69), .B(n67), .Y(SUM[22]) );
  AOI21X1 U72 ( .A(n145), .B(n70), .C(n71), .Y(n67) );
  NAND2X1 U73 ( .A(n144), .B(n68), .Y(n69) );
  NAND2X1 U74 ( .A(B[22]), .B(A[22]), .Y(n68) );
  NOR2X1 U75 ( .A(B[22]), .B(A[22]), .Y(n66) );
  XOR2X1 U76 ( .A(n70), .B(n73), .Y(SUM[21]) );
  NOR2X1 U77 ( .A(n71), .B(n72), .Y(n73) );
  NOR2X1 U78 ( .A(B[21]), .B(A[21]), .Y(n72) );
  AND2X1 U79 ( .A(B[21]), .B(A[21]), .Y(n71) );
  OAI21X1 U80 ( .A(n74), .B(n75), .C(n76), .Y(n70) );
  XOR2X1 U81 ( .A(n77), .B(n75), .Y(SUM[20]) );
  AOI21X1 U82 ( .A(n147), .B(n78), .C(n79), .Y(n75) );
  NAND2X1 U83 ( .A(n146), .B(n76), .Y(n77) );
  NAND2X1 U84 ( .A(B[20]), .B(A[20]), .Y(n76) );
  NOR2X1 U85 ( .A(B[20]), .B(A[20]), .Y(n74) );
  XOR2X1 U86 ( .A(n78), .B(n81), .Y(SUM[19]) );
  NOR2X1 U87 ( .A(n79), .B(n80), .Y(n81) );
  NOR2X1 U88 ( .A(B[19]), .B(A[19]), .Y(n80) );
  AND2X1 U89 ( .A(B[19]), .B(A[19]), .Y(n79) );
  OAI21X1 U90 ( .A(n82), .B(n83), .C(n84), .Y(n78) );
  XOR2X1 U91 ( .A(n85), .B(n83), .Y(SUM[18]) );
  AOI21X1 U92 ( .A(n149), .B(n86), .C(n87), .Y(n83) );
  NAND2X1 U93 ( .A(n148), .B(n84), .Y(n85) );
  NAND2X1 U94 ( .A(B[18]), .B(A[18]), .Y(n84) );
  NOR2X1 U95 ( .A(B[18]), .B(A[18]), .Y(n82) );
  XOR2X1 U96 ( .A(n86), .B(n89), .Y(SUM[17]) );
  NOR2X1 U97 ( .A(n87), .B(n88), .Y(n89) );
  NOR2X1 U98 ( .A(B[17]), .B(A[17]), .Y(n88) );
  AND2X1 U99 ( .A(B[17]), .B(A[17]), .Y(n87) );
  OAI21X1 U100 ( .A(n90), .B(n91), .C(n92), .Y(n86) );
  XOR2X1 U101 ( .A(n93), .B(n91), .Y(SUM[16]) );
  AOI21X1 U102 ( .A(n122), .B(n94), .C(n95), .Y(n91) );
  NAND2X1 U103 ( .A(n121), .B(n92), .Y(n93) );
  NAND2X1 U104 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NOR2X1 U105 ( .A(B[16]), .B(A[16]), .Y(n90) );
  XOR2X1 U106 ( .A(n94), .B(n97), .Y(SUM[15]) );
  NOR2X1 U107 ( .A(n95), .B(n96), .Y(n97) );
  NOR2X1 U108 ( .A(B[15]), .B(A[15]), .Y(n96) );
  AND2X1 U109 ( .A(B[15]), .B(A[15]), .Y(n95) );
  OAI21X1 U110 ( .A(n98), .B(n99), .C(n100), .Y(n94) );
  XOR2X1 U111 ( .A(n101), .B(n99), .Y(SUM[14]) );
  AOI21X1 U112 ( .A(n124), .B(n102), .C(n103), .Y(n99) );
  NAND2X1 U113 ( .A(n123), .B(n100), .Y(n101) );
  NAND2X1 U114 ( .A(B[14]), .B(A[14]), .Y(n100) );
  NOR2X1 U115 ( .A(B[14]), .B(A[14]), .Y(n98) );
  XOR2X1 U116 ( .A(n102), .B(n105), .Y(SUM[13]) );
  NOR2X1 U117 ( .A(n103), .B(n104), .Y(n105) );
  NOR2X1 U118 ( .A(B[13]), .B(A[13]), .Y(n104) );
  AND2X1 U119 ( .A(B[13]), .B(A[13]), .Y(n103) );
  OAI21X1 U120 ( .A(n106), .B(n126), .C(n107), .Y(n102) );
  XOR2X1 U121 ( .A(n108), .B(n126), .Y(SUM[12]) );
  OAI21X1 U122 ( .A(n110), .B(n111), .C(n112), .Y(n109) );
  AOI21X1 U123 ( .A(n113), .B(n129), .C(n128), .Y(n111) );
  NAND2X1 U124 ( .A(n125), .B(n107), .Y(n108) );
  NAND2X1 U125 ( .A(B[12]), .B(A[12]), .Y(n107) );
  NOR2X1 U126 ( .A(B[12]), .B(A[12]), .Y(n106) );
  XOR2X1 U127 ( .A(n115), .B(n116), .Y(SUM[11]) );
  NOR2X1 U128 ( .A(n127), .B(n110), .Y(n116) );
  NOR2X1 U129 ( .A(B[11]), .B(A[11]), .Y(n110) );
  NAND2X1 U130 ( .A(B[11]), .B(A[11]), .Y(n112) );
  OAI21X1 U131 ( .A(n117), .B(n131), .C(n114), .Y(n115) );
  XOR2X1 U132 ( .A(n118), .B(n131), .Y(SUM[10]) );
  OAI21X1 U133 ( .A(n132), .B(n32), .C(n33), .Y(n113) );
  NAND2X1 U134 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NOR2X1 U135 ( .A(B[9]), .B(A[9]), .Y(n32) );
  OAI21X1 U136 ( .A(n36), .B(n134), .C(n35), .Y(n30) );
  NAND2X1 U137 ( .A(B[8]), .B(A[8]), .Y(n35) );
  OAI21X1 U138 ( .A(n37), .B(n135), .C(n120), .Y(n119) );
  OAI21X1 U139 ( .A(n141), .B(A[7]), .C(B[7]), .Y(n120) );
  NAND2X1 U140 ( .A(B[6]), .B(A[6]), .Y(n37) );
  NOR2X1 U141 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NAND2X1 U142 ( .A(n129), .B(n114), .Y(n118) );
  NAND2X1 U143 ( .A(B[10]), .B(A[10]), .Y(n114) );
  NOR2X1 U144 ( .A(B[10]), .B(A[10]), .Y(n117) );
  INVX2 U2 ( .A(n90), .Y(n121) );
  INVX2 U3 ( .A(n96), .Y(n122) );
  INVX2 U4 ( .A(n98), .Y(n123) );
  INVX2 U5 ( .A(n104), .Y(n124) );
  INVX2 U6 ( .A(n106), .Y(n125) );
  INVX2 U7 ( .A(n109), .Y(n126) );
  INVX2 U8 ( .A(n112), .Y(n127) );
  INVX2 U9 ( .A(n114), .Y(n128) );
  INVX2 U10 ( .A(n117), .Y(n129) );
  INVX2 U11 ( .A(n33), .Y(n130) );
  INVX2 U12 ( .A(n113), .Y(n131) );
  INVX2 U13 ( .A(n30), .Y(n132) );
  INVX2 U14 ( .A(n36), .Y(n133) );
  INVX2 U15 ( .A(n119), .Y(n134) );
  INVX2 U16 ( .A(A[7]), .Y(n135) );
  INVX2 U17 ( .A(n42), .Y(n136) );
  INVX2 U18 ( .A(n48), .Y(n137) );
  INVX2 U19 ( .A(n50), .Y(n138) );
  INVX2 U20 ( .A(n56), .Y(n139) );
  INVX2 U21 ( .A(n39), .Y(SUM[6]) );
  INVX2 U22 ( .A(n37), .Y(n141) );
  INVX2 U23 ( .A(n58), .Y(n142) );
  INVX2 U24 ( .A(n64), .Y(n143) );
  INVX2 U25 ( .A(n66), .Y(n144) );
  INVX2 U26 ( .A(n72), .Y(n145) );
  INVX2 U27 ( .A(n74), .Y(n146) );
  INVX2 U28 ( .A(n80), .Y(n147) );
  INVX2 U29 ( .A(n82), .Y(n148) );
  INVX2 U30 ( .A(n88), .Y(n149) );
endmodule


module CannyEdge_DW02_mult_20 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] , \ab[7][27] ,
         \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][31] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][31] , \ab[3][30] ,
         \ab[3][29] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] , \ab[2][27] ,
         \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][31] ,
         \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] ,
         \ab[0][25] , \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] ,
         \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] ,
         \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] ,
         \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] ,
         \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] ,
         \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[30] , n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n110, n111, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S14_31_0 ( .A(n117), .B(\CARRYB[7][23] ), .C(\SUMB[7][24] ), .YC(
        \A2[30] ), .YS(\A1[29] ) );
  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S4_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S4_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S4_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S4_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  FAX1 S4_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S4_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S4_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S4_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  FAX1 S4_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S4_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S4_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S4_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  FAX1 S4_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S4_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S4_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S4_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  FAX1 S4_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S4_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S4_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S4_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  FAX1 S4_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S4_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S5_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .C(\ab[6][31] ), .YC(
        \CARRYB[7][30] ), .YS(\SUMB[7][30] ) );
  FAX1 S14_31 ( .A(QA), .B(QB), .C(\ab[7][31] ), .YC(\CARRYB[7][31] ), .YS(
        \SUMB[7][31] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  FAX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  FAX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  FAX1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  FAX1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  FAX1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .C(\ab[5][31] ), .YC(
        \CARRYB[6][30] ), .YS(\SUMB[6][30] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .C(\ab[4][31] ), .YC(
        \CARRYB[5][30] ), .YS(\SUMB[5][30] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .C(\ab[3][31] ), .YC(
        \CARRYB[4][30] ), .YS(\SUMB[4][30] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .C(\ab[2][31] ), .YC(
        \CARRYB[3][30] ), .YS(\SUMB[3][30] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n42), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n41), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n40), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n39), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n38), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n37), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n36), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n35), .C(\SUMB[1][8] ), .YC(\CARRYB[2][7] ), 
        .YS(\SUMB[2][7] ) );
  FAX1 S2_2_8 ( .A(\ab[2][8] ), .B(n34), .C(\SUMB[1][9] ), .YC(\CARRYB[2][8] ), 
        .YS(\SUMB[2][8] ) );
  FAX1 S2_2_9 ( .A(\ab[2][9] ), .B(n33), .C(\SUMB[1][10] ), .YC(\CARRYB[2][9] ), .YS(\SUMB[2][9] ) );
  FAX1 S2_2_10 ( .A(\ab[2][10] ), .B(n32), .C(\SUMB[1][11] ), .YC(
        \CARRYB[2][10] ), .YS(\SUMB[2][10] ) );
  FAX1 S2_2_11 ( .A(\ab[2][11] ), .B(n31), .C(\SUMB[1][12] ), .YC(
        \CARRYB[2][11] ), .YS(\SUMB[2][11] ) );
  FAX1 S2_2_12 ( .A(\ab[2][12] ), .B(n30), .C(\SUMB[1][13] ), .YC(
        \CARRYB[2][12] ), .YS(\SUMB[2][12] ) );
  FAX1 S2_2_13 ( .A(\ab[2][13] ), .B(n29), .C(\SUMB[1][14] ), .YC(
        \CARRYB[2][13] ), .YS(\SUMB[2][13] ) );
  FAX1 S2_2_14 ( .A(\ab[2][14] ), .B(n28), .C(\SUMB[1][15] ), .YC(
        \CARRYB[2][14] ), .YS(\SUMB[2][14] ) );
  FAX1 S2_2_15 ( .A(\ab[2][15] ), .B(n27), .C(\SUMB[1][16] ), .YC(
        \CARRYB[2][15] ), .YS(\SUMB[2][15] ) );
  FAX1 S2_2_16 ( .A(\ab[2][16] ), .B(n26), .C(\SUMB[1][17] ), .YC(
        \CARRYB[2][16] ), .YS(\SUMB[2][16] ) );
  FAX1 S2_2_17 ( .A(\ab[2][17] ), .B(n25), .C(\SUMB[1][18] ), .YC(
        \CARRYB[2][17] ), .YS(\SUMB[2][17] ) );
  FAX1 S2_2_18 ( .A(\ab[2][18] ), .B(n24), .C(\SUMB[1][19] ), .YC(
        \CARRYB[2][18] ), .YS(\SUMB[2][18] ) );
  FAX1 S2_2_19 ( .A(\ab[2][19] ), .B(n23), .C(\SUMB[1][20] ), .YC(
        \CARRYB[2][19] ), .YS(\SUMB[2][19] ) );
  FAX1 S2_2_20 ( .A(\ab[2][20] ), .B(n22), .C(\SUMB[1][21] ), .YC(
        \CARRYB[2][20] ), .YS(\SUMB[2][20] ) );
  FAX1 S2_2_21 ( .A(\ab[2][21] ), .B(n21), .C(\SUMB[1][22] ), .YC(
        \CARRYB[2][21] ), .YS(\SUMB[2][21] ) );
  FAX1 S2_2_22 ( .A(\ab[2][22] ), .B(n20), .C(\SUMB[1][23] ), .YC(
        \CARRYB[2][22] ), .YS(\SUMB[2][22] ) );
  FAX1 S2_2_23 ( .A(\ab[2][23] ), .B(n19), .C(\SUMB[1][24] ), .YC(
        \CARRYB[2][23] ), .YS(\SUMB[2][23] ) );
  FAX1 S2_2_24 ( .A(\ab[2][24] ), .B(n18), .C(\SUMB[1][25] ), .YC(
        \CARRYB[2][24] ), .YS(\SUMB[2][24] ) );
  FAX1 S2_2_25 ( .A(\ab[2][25] ), .B(n17), .C(\SUMB[1][26] ), .YC(
        \CARRYB[2][25] ), .YS(\SUMB[2][25] ) );
  FAX1 S2_2_26 ( .A(\ab[2][26] ), .B(n16), .C(\SUMB[1][27] ), .YC(
        \CARRYB[2][26] ), .YS(\SUMB[2][26] ) );
  FAX1 S2_2_27 ( .A(\ab[2][27] ), .B(n15), .C(\SUMB[1][28] ), .YC(
        \CARRYB[2][27] ), .YS(\SUMB[2][27] ) );
  FAX1 S2_2_28 ( .A(\ab[2][28] ), .B(n14), .C(\SUMB[1][29] ), .YC(
        \CARRYB[2][28] ), .YS(\SUMB[2][28] ) );
  FAX1 S2_2_29 ( .A(\ab[2][29] ), .B(n13), .C(\SUMB[1][30] ), .YC(
        \CARRYB[2][29] ), .YS(\SUMB[2][29] ) );
  FAX1 S3_2_30 ( .A(\ab[2][30] ), .B(n12), .C(\ab[1][31] ), .YC(
        \CARRYB[2][30] ), .YS(\SUMB[2][30] ) );
  AND2X2 U2 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(n3) );
  AND2X2 U3 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(n4) );
  AND2X2 U4 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(n5) );
  AND2X2 U5 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(n6) );
  AND2X2 U6 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(n7) );
  AND2X2 U7 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(n8) );
  AND2X2 U8 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(n9) );
  AND2X2 U9 ( .A(TC), .B(A[7]), .Y(n10) );
  AND2X2 U10 ( .A(A[7]), .B(n115), .Y(n11) );
  AND2X2 U11 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Y(n12) );
  AND2X2 U12 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Y(n13) );
  AND2X2 U13 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Y(n24) );
  AND2X2 U24 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Y(n25) );
  AND2X2 U25 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Y(n26) );
  AND2X2 U26 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Y(n27) );
  AND2X2 U27 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n28) );
  AND2X2 U28 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n29) );
  AND2X2 U29 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n30) );
  AND2X2 U30 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Y(n31) );
  AND2X2 U31 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n36) );
  AND2X2 U36 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n37) );
  AND2X2 U37 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n38) );
  AND2X2 U38 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n39) );
  AND2X2 U39 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n40) );
  AND2X2 U40 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n41) );
  AND2X2 U41 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n42) );
  AND2X2 U42 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][0] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(n53) );
  AND2X2 U53 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(n54) );
  AND2X2 U54 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(n55) );
  AND2X2 U55 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(n56) );
  AND2X2 U56 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(n57) );
  AND2X2 U57 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(n58) );
  AND2X2 U58 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(n59) );
  AND2X2 U59 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(n60) );
  AND2X2 U60 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(n61) );
  AND2X2 U61 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(n62) );
  AND2X2 U62 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(n63) );
  AND2X2 U63 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n64) );
  AND2X2 U64 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(n65) );
  AND2X2 U65 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(n66) );
  XOR2X1 U68 ( .A(\SUMB[7][0] ), .B(n10), .Y(\A1[5] ) );
  XOR2X1 U69 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  XOR2X1 U70 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  XOR2X1 U71 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  XOR2X1 U72 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  XOR2X1 U73 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  XOR2X1 U74 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  XOR2X1 U75 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  XOR2X1 U76 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  XOR2X1 U77 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  XOR2X1 U78 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  XOR2X1 U79 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  XOR2X1 U80 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  XOR2X1 U81 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  XOR2X1 U82 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  XOR2X1 U83 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  XOR2X1 U84 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  XOR2X1 U85 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  XOR2X1 U86 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  XOR2X1 U87 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  XOR2X1 U88 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  XOR2X1 U89 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  XOR2X1 U90 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  XOR2X1 U91 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  XOR2X1 U92 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  XOR2X1 U93 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  XOR2X1 U94 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  XOR2X1 U95 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  XOR2X1 U96 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  XOR2X1 U97 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  XOR2X1 U98 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(\A1[36] ) );
  XOR2X1 U99 ( .A(\CARRYB[7][31] ), .B(TC), .Y(\A1[37] ) );
  XOR2X1 U100 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U101 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U102 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U103 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U104 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U105 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U106 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U107 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  XOR2X1 U108 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(\SUMB[1][8] ) );
  XOR2X1 U109 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Y(\SUMB[1][9] ) );
  XOR2X1 U110 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Y(\SUMB[1][10] ) );
  XOR2X1 U111 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U112 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Y(\SUMB[1][12] ) );
  XOR2X1 U113 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  XOR2X1 U114 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  XOR2X1 U115 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Y(\SUMB[1][15] ) );
  XOR2X1 U116 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Y(\SUMB[1][16] ) );
  XOR2X1 U117 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Y(\SUMB[1][17] ) );
  XOR2X1 U118 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Y(\SUMB[1][18] ) );
  XOR2X1 U119 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Y(\SUMB[1][19] ) );
  XOR2X1 U120 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Y(\SUMB[1][20] ) );
  XOR2X1 U121 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Y(\SUMB[1][21] ) );
  XOR2X1 U122 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Y(\SUMB[1][22] ) );
  XOR2X1 U123 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Y(\SUMB[1][23] ) );
  XOR2X1 U124 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Y(\SUMB[1][24] ) );
  XOR2X1 U125 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Y(\SUMB[1][25] ) );
  XOR2X1 U126 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Y(\SUMB[1][26] ) );
  XOR2X1 U127 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Y(\SUMB[1][27] ) );
  XOR2X1 U128 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Y(\SUMB[1][28] ) );
  XOR2X1 U129 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Y(\SUMB[1][29] ) );
  XOR2X1 U130 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Y(\SUMB[1][30] ) );
  MUX2X1 U171 ( .B(n116), .A(n114), .S(B[9]), .Y(\ab[7][9] ) );
  MUX2X1 U172 ( .B(n116), .A(n114), .S(B[8]), .Y(\ab[7][8] ) );
  MUX2X1 U173 ( .B(n116), .A(n114), .S(B[7]), .Y(\ab[7][7] ) );
  MUX2X1 U174 ( .B(n116), .A(n114), .S(B[6]), .Y(\ab[7][6] ) );
  MUX2X1 U175 ( .B(n116), .A(n114), .S(B[5]), .Y(\ab[7][5] ) );
  MUX2X1 U176 ( .B(n116), .A(n114), .S(B[4]), .Y(\ab[7][4] ) );
  MUX2X1 U177 ( .B(n116), .A(n114), .S(B[3]), .Y(\ab[7][3] ) );
  AND2X1 U178 ( .A(A[7]), .B(B[31]), .Y(\ab[7][31] ) );
  MUX2X1 U179 ( .B(n116), .A(n114), .S(B[30]), .Y(\ab[7][30] ) );
  MUX2X1 U180 ( .B(n116), .A(n114), .S(B[2]), .Y(\ab[7][2] ) );
  MUX2X1 U181 ( .B(n116), .A(n114), .S(B[29]), .Y(\ab[7][29] ) );
  MUX2X1 U182 ( .B(n116), .A(n114), .S(B[28]), .Y(\ab[7][28] ) );
  MUX2X1 U183 ( .B(n116), .A(n114), .S(B[27]), .Y(\ab[7][27] ) );
  MUX2X1 U184 ( .B(n116), .A(n114), .S(B[26]), .Y(\ab[7][26] ) );
  MUX2X1 U185 ( .B(n116), .A(n114), .S(B[25]), .Y(\ab[7][25] ) );
  MUX2X1 U186 ( .B(n116), .A(n114), .S(B[24]), .Y(\ab[7][24] ) );
  MUX2X1 U187 ( .B(n116), .A(n114), .S(B[23]), .Y(\ab[7][23] ) );
  MUX2X1 U188 ( .B(n116), .A(n114), .S(B[22]), .Y(\ab[7][22] ) );
  MUX2X1 U189 ( .B(n116), .A(n114), .S(B[21]), .Y(\ab[7][21] ) );
  MUX2X1 U190 ( .B(n116), .A(n114), .S(B[20]), .Y(\ab[7][20] ) );
  MUX2X1 U191 ( .B(n116), .A(n114), .S(B[1]), .Y(\ab[7][1] ) );
  MUX2X1 U192 ( .B(n116), .A(n114), .S(B[19]), .Y(\ab[7][19] ) );
  MUX2X1 U193 ( .B(n116), .A(n114), .S(B[18]), .Y(\ab[7][18] ) );
  MUX2X1 U194 ( .B(n116), .A(n114), .S(B[17]), .Y(\ab[7][17] ) );
  MUX2X1 U195 ( .B(n116), .A(n114), .S(B[16]), .Y(\ab[7][16] ) );
  MUX2X1 U196 ( .B(n116), .A(n114), .S(B[15]), .Y(\ab[7][15] ) );
  MUX2X1 U197 ( .B(n116), .A(n114), .S(B[14]), .Y(\ab[7][14] ) );
  MUX2X1 U198 ( .B(n116), .A(n114), .S(B[13]), .Y(\ab[7][13] ) );
  MUX2X1 U199 ( .B(n116), .A(n114), .S(B[12]), .Y(\ab[7][12] ) );
  MUX2X1 U200 ( .B(n116), .A(n114), .S(B[11]), .Y(\ab[7][11] ) );
  MUX2X1 U201 ( .B(n116), .A(n114), .S(B[10]), .Y(\ab[7][10] ) );
  MUX2X1 U202 ( .B(n116), .A(n114), .S(B[0]), .Y(\ab[7][0] ) );
  NOR2X1 U203 ( .A(n147), .B(n155), .Y(\ab[6][9] ) );
  NOR2X1 U204 ( .A(n150), .B(n155), .Y(\ab[6][8] ) );
  NOR2X1 U205 ( .A(n118), .B(n155), .Y(\ab[6][7] ) );
  NOR2X1 U206 ( .A(n119), .B(n155), .Y(\ab[6][6] ) );
  NOR2X1 U207 ( .A(n120), .B(n155), .Y(\ab[6][5] ) );
  NOR2X1 U208 ( .A(n121), .B(n155), .Y(\ab[6][4] ) );
  NOR2X1 U209 ( .A(n122), .B(n155), .Y(\ab[6][3] ) );
  MUX2X1 U210 ( .B(n110), .A(n111), .S(A[6]), .Y(\ab[6][31] ) );
  NOR2X1 U211 ( .A(n146), .B(n155), .Y(\ab[6][30] ) );
  NOR2X1 U212 ( .A(n123), .B(n155), .Y(\ab[6][2] ) );
  NOR2X1 U213 ( .A(n145), .B(n155), .Y(\ab[6][29] ) );
  NOR2X1 U214 ( .A(n144), .B(n155), .Y(\ab[6][28] ) );
  NOR2X1 U215 ( .A(n143), .B(n155), .Y(\ab[6][27] ) );
  NOR2X1 U216 ( .A(n142), .B(n155), .Y(\ab[6][26] ) );
  NOR2X1 U217 ( .A(n141), .B(n155), .Y(\ab[6][25] ) );
  NOR2X1 U218 ( .A(n140), .B(n155), .Y(\ab[6][24] ) );
  NOR2X1 U219 ( .A(n139), .B(n155), .Y(\ab[6][23] ) );
  NOR2X1 U220 ( .A(n138), .B(n155), .Y(\ab[6][22] ) );
  NOR2X1 U221 ( .A(n137), .B(n155), .Y(\ab[6][21] ) );
  NOR2X1 U222 ( .A(n136), .B(n155), .Y(\ab[6][20] ) );
  NOR2X1 U223 ( .A(n124), .B(n155), .Y(\ab[6][1] ) );
  NOR2X1 U224 ( .A(n135), .B(n155), .Y(\ab[6][19] ) );
  NOR2X1 U225 ( .A(n134), .B(n155), .Y(\ab[6][18] ) );
  NOR2X1 U226 ( .A(n133), .B(n155), .Y(\ab[6][17] ) );
  NOR2X1 U227 ( .A(n132), .B(n155), .Y(\ab[6][16] ) );
  NOR2X1 U228 ( .A(n131), .B(n155), .Y(\ab[6][15] ) );
  NOR2X1 U229 ( .A(n130), .B(n155), .Y(\ab[6][14] ) );
  NOR2X1 U230 ( .A(n129), .B(n155), .Y(\ab[6][13] ) );
  NOR2X1 U231 ( .A(n128), .B(n155), .Y(\ab[6][12] ) );
  NOR2X1 U232 ( .A(n127), .B(n155), .Y(\ab[6][11] ) );
  NOR2X1 U233 ( .A(n148), .B(n155), .Y(\ab[6][10] ) );
  NOR2X1 U234 ( .A(n125), .B(n155), .Y(\ab[6][0] ) );
  NOR2X1 U235 ( .A(n147), .B(n154), .Y(\ab[5][9] ) );
  NOR2X1 U236 ( .A(n150), .B(n154), .Y(\ab[5][8] ) );
  NOR2X1 U237 ( .A(n118), .B(n154), .Y(\ab[5][7] ) );
  NOR2X1 U238 ( .A(n119), .B(n154), .Y(\ab[5][6] ) );
  NOR2X1 U239 ( .A(n120), .B(n154), .Y(\ab[5][5] ) );
  NOR2X1 U240 ( .A(n121), .B(n154), .Y(\ab[5][4] ) );
  NOR2X1 U241 ( .A(n122), .B(n154), .Y(\ab[5][3] ) );
  MUX2X1 U242 ( .B(n110), .A(n111), .S(A[5]), .Y(\ab[5][31] ) );
  NOR2X1 U243 ( .A(n146), .B(n154), .Y(\ab[5][30] ) );
  NOR2X1 U244 ( .A(n123), .B(n154), .Y(\ab[5][2] ) );
  NOR2X1 U245 ( .A(n145), .B(n154), .Y(\ab[5][29] ) );
  NOR2X1 U246 ( .A(n144), .B(n154), .Y(\ab[5][28] ) );
  NOR2X1 U247 ( .A(n143), .B(n154), .Y(\ab[5][27] ) );
  NOR2X1 U248 ( .A(n142), .B(n154), .Y(\ab[5][26] ) );
  NOR2X1 U249 ( .A(n141), .B(n154), .Y(\ab[5][25] ) );
  NOR2X1 U250 ( .A(n140), .B(n154), .Y(\ab[5][24] ) );
  NOR2X1 U251 ( .A(n139), .B(n154), .Y(\ab[5][23] ) );
  NOR2X1 U252 ( .A(n138), .B(n154), .Y(\ab[5][22] ) );
  NOR2X1 U253 ( .A(n137), .B(n154), .Y(\ab[5][21] ) );
  NOR2X1 U254 ( .A(n136), .B(n154), .Y(\ab[5][20] ) );
  NOR2X1 U255 ( .A(n124), .B(n154), .Y(\ab[5][1] ) );
  NOR2X1 U256 ( .A(n135), .B(n154), .Y(\ab[5][19] ) );
  NOR2X1 U257 ( .A(n134), .B(n154), .Y(\ab[5][18] ) );
  NOR2X1 U258 ( .A(n133), .B(n154), .Y(\ab[5][17] ) );
  NOR2X1 U259 ( .A(n132), .B(n154), .Y(\ab[5][16] ) );
  NOR2X1 U260 ( .A(n131), .B(n154), .Y(\ab[5][15] ) );
  NOR2X1 U261 ( .A(n130), .B(n154), .Y(\ab[5][14] ) );
  NOR2X1 U262 ( .A(n129), .B(n154), .Y(\ab[5][13] ) );
  NOR2X1 U263 ( .A(n128), .B(n154), .Y(\ab[5][12] ) );
  NOR2X1 U264 ( .A(n127), .B(n154), .Y(\ab[5][11] ) );
  NOR2X1 U265 ( .A(n148), .B(n154), .Y(\ab[5][10] ) );
  NOR2X1 U266 ( .A(n125), .B(n154), .Y(\ab[5][0] ) );
  NOR2X1 U267 ( .A(n147), .B(n153), .Y(\ab[4][9] ) );
  NOR2X1 U268 ( .A(n150), .B(n153), .Y(\ab[4][8] ) );
  NOR2X1 U269 ( .A(n118), .B(n153), .Y(\ab[4][7] ) );
  NOR2X1 U270 ( .A(n119), .B(n153), .Y(\ab[4][6] ) );
  NOR2X1 U271 ( .A(n120), .B(n153), .Y(\ab[4][5] ) );
  NOR2X1 U272 ( .A(n121), .B(n153), .Y(\ab[4][4] ) );
  NOR2X1 U273 ( .A(n122), .B(n153), .Y(\ab[4][3] ) );
  MUX2X1 U274 ( .B(n110), .A(n111), .S(A[4]), .Y(\ab[4][31] ) );
  NOR2X1 U275 ( .A(n146), .B(n153), .Y(\ab[4][30] ) );
  NOR2X1 U276 ( .A(n123), .B(n153), .Y(\ab[4][2] ) );
  NOR2X1 U277 ( .A(n145), .B(n153), .Y(\ab[4][29] ) );
  NOR2X1 U278 ( .A(n144), .B(n153), .Y(\ab[4][28] ) );
  NOR2X1 U279 ( .A(n143), .B(n153), .Y(\ab[4][27] ) );
  NOR2X1 U280 ( .A(n142), .B(n153), .Y(\ab[4][26] ) );
  NOR2X1 U281 ( .A(n141), .B(n153), .Y(\ab[4][25] ) );
  NOR2X1 U282 ( .A(n140), .B(n153), .Y(\ab[4][24] ) );
  NOR2X1 U283 ( .A(n139), .B(n153), .Y(\ab[4][23] ) );
  NOR2X1 U284 ( .A(n138), .B(n153), .Y(\ab[4][22] ) );
  NOR2X1 U285 ( .A(n137), .B(n153), .Y(\ab[4][21] ) );
  NOR2X1 U286 ( .A(n136), .B(n153), .Y(\ab[4][20] ) );
  NOR2X1 U287 ( .A(n124), .B(n153), .Y(\ab[4][1] ) );
  NOR2X1 U288 ( .A(n135), .B(n153), .Y(\ab[4][19] ) );
  NOR2X1 U289 ( .A(n134), .B(n153), .Y(\ab[4][18] ) );
  NOR2X1 U290 ( .A(n133), .B(n153), .Y(\ab[4][17] ) );
  NOR2X1 U291 ( .A(n132), .B(n153), .Y(\ab[4][16] ) );
  NOR2X1 U292 ( .A(n131), .B(n153), .Y(\ab[4][15] ) );
  NOR2X1 U293 ( .A(n130), .B(n153), .Y(\ab[4][14] ) );
  NOR2X1 U294 ( .A(n129), .B(n153), .Y(\ab[4][13] ) );
  NOR2X1 U295 ( .A(n128), .B(n153), .Y(\ab[4][12] ) );
  NOR2X1 U296 ( .A(n127), .B(n153), .Y(\ab[4][11] ) );
  NOR2X1 U297 ( .A(n148), .B(n153), .Y(\ab[4][10] ) );
  NOR2X1 U298 ( .A(n125), .B(n153), .Y(\ab[4][0] ) );
  NOR2X1 U299 ( .A(n147), .B(n152), .Y(\ab[3][9] ) );
  NOR2X1 U300 ( .A(n150), .B(n152), .Y(\ab[3][8] ) );
  NOR2X1 U301 ( .A(n118), .B(n152), .Y(\ab[3][7] ) );
  NOR2X1 U302 ( .A(n119), .B(n152), .Y(\ab[3][6] ) );
  NOR2X1 U303 ( .A(n120), .B(n152), .Y(\ab[3][5] ) );
  NOR2X1 U304 ( .A(n121), .B(n152), .Y(\ab[3][4] ) );
  NOR2X1 U305 ( .A(n122), .B(n152), .Y(\ab[3][3] ) );
  MUX2X1 U306 ( .B(n110), .A(n111), .S(A[3]), .Y(\ab[3][31] ) );
  NOR2X1 U307 ( .A(n146), .B(n152), .Y(\ab[3][30] ) );
  NOR2X1 U308 ( .A(n123), .B(n152), .Y(\ab[3][2] ) );
  NOR2X1 U309 ( .A(n145), .B(n152), .Y(\ab[3][29] ) );
  NOR2X1 U310 ( .A(n144), .B(n152), .Y(\ab[3][28] ) );
  NOR2X1 U311 ( .A(n143), .B(n152), .Y(\ab[3][27] ) );
  NOR2X1 U312 ( .A(n142), .B(n152), .Y(\ab[3][26] ) );
  NOR2X1 U313 ( .A(n141), .B(n152), .Y(\ab[3][25] ) );
  NOR2X1 U314 ( .A(n140), .B(n152), .Y(\ab[3][24] ) );
  NOR2X1 U315 ( .A(n139), .B(n152), .Y(\ab[3][23] ) );
  NOR2X1 U316 ( .A(n138), .B(n152), .Y(\ab[3][22] ) );
  NOR2X1 U317 ( .A(n137), .B(n152), .Y(\ab[3][21] ) );
  NOR2X1 U318 ( .A(n136), .B(n152), .Y(\ab[3][20] ) );
  NOR2X1 U319 ( .A(n124), .B(n152), .Y(\ab[3][1] ) );
  NOR2X1 U320 ( .A(n135), .B(n152), .Y(\ab[3][19] ) );
  NOR2X1 U321 ( .A(n134), .B(n152), .Y(\ab[3][18] ) );
  NOR2X1 U322 ( .A(n133), .B(n152), .Y(\ab[3][17] ) );
  NOR2X1 U323 ( .A(n132), .B(n152), .Y(\ab[3][16] ) );
  NOR2X1 U324 ( .A(n131), .B(n152), .Y(\ab[3][15] ) );
  NOR2X1 U325 ( .A(n130), .B(n152), .Y(\ab[3][14] ) );
  NOR2X1 U326 ( .A(n129), .B(n152), .Y(\ab[3][13] ) );
  NOR2X1 U327 ( .A(n128), .B(n152), .Y(\ab[3][12] ) );
  NOR2X1 U328 ( .A(n127), .B(n152), .Y(\ab[3][11] ) );
  NOR2X1 U329 ( .A(n148), .B(n152), .Y(\ab[3][10] ) );
  NOR2X1 U330 ( .A(n125), .B(n152), .Y(\ab[3][0] ) );
  NOR2X1 U331 ( .A(n147), .B(n149), .Y(\ab[2][9] ) );
  NOR2X1 U332 ( .A(n150), .B(n149), .Y(\ab[2][8] ) );
  NOR2X1 U333 ( .A(n118), .B(n149), .Y(\ab[2][7] ) );
  NOR2X1 U334 ( .A(n119), .B(n149), .Y(\ab[2][6] ) );
  NOR2X1 U335 ( .A(n120), .B(n149), .Y(\ab[2][5] ) );
  NOR2X1 U336 ( .A(n121), .B(n149), .Y(\ab[2][4] ) );
  NOR2X1 U337 ( .A(n122), .B(n149), .Y(\ab[2][3] ) );
  MUX2X1 U338 ( .B(n110), .A(n111), .S(A[2]), .Y(\ab[2][31] ) );
  NOR2X1 U339 ( .A(n146), .B(n149), .Y(\ab[2][30] ) );
  NOR2X1 U340 ( .A(n123), .B(n149), .Y(\ab[2][2] ) );
  NOR2X1 U341 ( .A(n145), .B(n149), .Y(\ab[2][29] ) );
  NOR2X1 U342 ( .A(n144), .B(n149), .Y(\ab[2][28] ) );
  NOR2X1 U343 ( .A(n143), .B(n149), .Y(\ab[2][27] ) );
  NOR2X1 U344 ( .A(n142), .B(n149), .Y(\ab[2][26] ) );
  NOR2X1 U345 ( .A(n141), .B(n149), .Y(\ab[2][25] ) );
  NOR2X1 U346 ( .A(n140), .B(n149), .Y(\ab[2][24] ) );
  NOR2X1 U347 ( .A(n139), .B(n149), .Y(\ab[2][23] ) );
  NOR2X1 U348 ( .A(n138), .B(n149), .Y(\ab[2][22] ) );
  NOR2X1 U349 ( .A(n137), .B(n149), .Y(\ab[2][21] ) );
  NOR2X1 U350 ( .A(n136), .B(n149), .Y(\ab[2][20] ) );
  NOR2X1 U351 ( .A(n124), .B(n149), .Y(\ab[2][1] ) );
  NOR2X1 U352 ( .A(n135), .B(n149), .Y(\ab[2][19] ) );
  NOR2X1 U353 ( .A(n134), .B(n149), .Y(\ab[2][18] ) );
  NOR2X1 U354 ( .A(n133), .B(n149), .Y(\ab[2][17] ) );
  NOR2X1 U355 ( .A(n132), .B(n149), .Y(\ab[2][16] ) );
  NOR2X1 U356 ( .A(n131), .B(n149), .Y(\ab[2][15] ) );
  NOR2X1 U357 ( .A(n130), .B(n149), .Y(\ab[2][14] ) );
  NOR2X1 U358 ( .A(n129), .B(n149), .Y(\ab[2][13] ) );
  NOR2X1 U359 ( .A(n128), .B(n149), .Y(\ab[2][12] ) );
  NOR2X1 U360 ( .A(n127), .B(n149), .Y(\ab[2][11] ) );
  NOR2X1 U361 ( .A(n148), .B(n149), .Y(\ab[2][10] ) );
  NOR2X1 U362 ( .A(n125), .B(n149), .Y(\ab[2][0] ) );
  NOR2X1 U363 ( .A(n147), .B(n151), .Y(\ab[1][9] ) );
  NOR2X1 U364 ( .A(n150), .B(n151), .Y(\ab[1][8] ) );
  NOR2X1 U365 ( .A(n118), .B(n151), .Y(\ab[1][7] ) );
  NOR2X1 U366 ( .A(n119), .B(n151), .Y(\ab[1][6] ) );
  NOR2X1 U367 ( .A(n120), .B(n151), .Y(\ab[1][5] ) );
  NOR2X1 U368 ( .A(n121), .B(n151), .Y(\ab[1][4] ) );
  NOR2X1 U369 ( .A(n122), .B(n151), .Y(\ab[1][3] ) );
  MUX2X1 U370 ( .B(n110), .A(n111), .S(A[1]), .Y(\ab[1][31] ) );
  NOR2X1 U371 ( .A(n146), .B(n151), .Y(\ab[1][30] ) );
  NOR2X1 U372 ( .A(n123), .B(n151), .Y(\ab[1][2] ) );
  NOR2X1 U373 ( .A(n145), .B(n151), .Y(\ab[1][29] ) );
  NOR2X1 U374 ( .A(n144), .B(n151), .Y(\ab[1][28] ) );
  NOR2X1 U375 ( .A(n143), .B(n151), .Y(\ab[1][27] ) );
  NOR2X1 U376 ( .A(n142), .B(n151), .Y(\ab[1][26] ) );
  NOR2X1 U377 ( .A(n141), .B(n151), .Y(\ab[1][25] ) );
  NOR2X1 U378 ( .A(n140), .B(n151), .Y(\ab[1][24] ) );
  NOR2X1 U379 ( .A(n139), .B(n151), .Y(\ab[1][23] ) );
  NOR2X1 U380 ( .A(n138), .B(n151), .Y(\ab[1][22] ) );
  NOR2X1 U381 ( .A(n137), .B(n151), .Y(\ab[1][21] ) );
  NOR2X1 U382 ( .A(n136), .B(n151), .Y(\ab[1][20] ) );
  NOR2X1 U383 ( .A(n124), .B(n151), .Y(\ab[1][1] ) );
  NOR2X1 U384 ( .A(n135), .B(n151), .Y(\ab[1][19] ) );
  NOR2X1 U385 ( .A(n134), .B(n151), .Y(\ab[1][18] ) );
  NOR2X1 U386 ( .A(n133), .B(n151), .Y(\ab[1][17] ) );
  NOR2X1 U387 ( .A(n132), .B(n151), .Y(\ab[1][16] ) );
  NOR2X1 U388 ( .A(n131), .B(n151), .Y(\ab[1][15] ) );
  NOR2X1 U389 ( .A(n130), .B(n151), .Y(\ab[1][14] ) );
  NOR2X1 U390 ( .A(n129), .B(n151), .Y(\ab[1][13] ) );
  NOR2X1 U391 ( .A(n128), .B(n151), .Y(\ab[1][12] ) );
  NOR2X1 U392 ( .A(n127), .B(n151), .Y(\ab[1][11] ) );
  NOR2X1 U393 ( .A(n148), .B(n151), .Y(\ab[1][10] ) );
  NOR2X1 U394 ( .A(n125), .B(n151), .Y(\ab[1][0] ) );
  NOR2X1 U395 ( .A(n147), .B(n126), .Y(\ab[0][9] ) );
  NOR2X1 U396 ( .A(n150), .B(n126), .Y(\ab[0][8] ) );
  NOR2X1 U397 ( .A(n118), .B(n126), .Y(\ab[0][7] ) );
  NOR2X1 U398 ( .A(n119), .B(n126), .Y(\ab[0][6] ) );
  NOR2X1 U399 ( .A(n120), .B(n126), .Y(\ab[0][5] ) );
  NOR2X1 U400 ( .A(n121), .B(n126), .Y(\ab[0][4] ) );
  NOR2X1 U401 ( .A(n122), .B(n126), .Y(\ab[0][3] ) );
  MUX2X1 U402 ( .B(n110), .A(n111), .S(A[0]), .Y(\ab[0][31] ) );
  NAND2X1 U403 ( .A(B[31]), .B(n115), .Y(n111) );
  NOR2X1 U404 ( .A(n146), .B(n126), .Y(\ab[0][30] ) );
  NOR2X1 U405 ( .A(n123), .B(n126), .Y(\ab[0][2] ) );
  NOR2X1 U406 ( .A(n145), .B(n126), .Y(\ab[0][29] ) );
  NOR2X1 U407 ( .A(n144), .B(n126), .Y(\ab[0][28] ) );
  NOR2X1 U408 ( .A(n143), .B(n126), .Y(\ab[0][27] ) );
  NOR2X1 U409 ( .A(n142), .B(n126), .Y(\ab[0][26] ) );
  NOR2X1 U410 ( .A(n141), .B(n126), .Y(\ab[0][25] ) );
  NOR2X1 U411 ( .A(n140), .B(n126), .Y(\ab[0][24] ) );
  NOR2X1 U412 ( .A(n139), .B(n126), .Y(\ab[0][23] ) );
  NOR2X1 U413 ( .A(n138), .B(n126), .Y(\ab[0][22] ) );
  NOR2X1 U414 ( .A(n137), .B(n126), .Y(\ab[0][21] ) );
  NOR2X1 U415 ( .A(n136), .B(n126), .Y(\ab[0][20] ) );
  NOR2X1 U416 ( .A(n124), .B(n126), .Y(\ab[0][1] ) );
  NOR2X1 U417 ( .A(n135), .B(n126), .Y(\ab[0][19] ) );
  NOR2X1 U418 ( .A(n134), .B(n126), .Y(\ab[0][18] ) );
  NOR2X1 U419 ( .A(n133), .B(n126), .Y(\ab[0][17] ) );
  NOR2X1 U420 ( .A(n132), .B(n126), .Y(\ab[0][16] ) );
  NOR2X1 U421 ( .A(n131), .B(n126), .Y(\ab[0][15] ) );
  NOR2X1 U422 ( .A(n130), .B(n126), .Y(\ab[0][14] ) );
  NOR2X1 U423 ( .A(n129), .B(n126), .Y(\ab[0][13] ) );
  NOR2X1 U424 ( .A(n128), .B(n126), .Y(\ab[0][12] ) );
  NOR2X1 U425 ( .A(n127), .B(n126), .Y(\ab[0][11] ) );
  NOR2X1 U426 ( .A(n148), .B(n126), .Y(\ab[0][10] ) );
  NAND2X1 U427 ( .A(B[31]), .B(TC), .Y(n110) );
  NOR2X1 U428 ( .A(B[31]), .B(n115), .Y(QB) );
  NOR2X1 U429 ( .A(A[7]), .B(n115), .Y(QA) );
  NOR2X1 U430 ( .A(n125), .B(n126), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_42 FS_1 ( .A({\A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n9, n8, n7, 
        n6, n5, n4, n3, \A2[30] , n45, n54, n46, n55, n47, n56, n48, n57, n49, 
        n58, n50, n59, n51, n60, n52, n61, n53, n62, n63, n66, n64, n65, n43, 
        n44, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  INVX2 U131 ( .A(n11), .Y(n114) );
  INVX2 U132 ( .A(TC), .Y(n115) );
  INVX2 U133 ( .A(n10), .Y(n116) );
  INVX2 U134 ( .A(n110), .Y(n117) );
  INVX2 U135 ( .A(B[7]), .Y(n118) );
  INVX2 U136 ( .A(B[6]), .Y(n119) );
  INVX2 U137 ( .A(B[5]), .Y(n120) );
  INVX2 U138 ( .A(B[4]), .Y(n121) );
  INVX2 U139 ( .A(B[3]), .Y(n122) );
  INVX2 U140 ( .A(B[2]), .Y(n123) );
  INVX2 U141 ( .A(B[1]), .Y(n124) );
  INVX2 U142 ( .A(B[0]), .Y(n125) );
  INVX2 U143 ( .A(A[0]), .Y(n126) );
  INVX2 U144 ( .A(B[11]), .Y(n127) );
  INVX2 U145 ( .A(B[12]), .Y(n128) );
  INVX2 U146 ( .A(B[13]), .Y(n129) );
  INVX2 U147 ( .A(B[14]), .Y(n130) );
  INVX2 U148 ( .A(B[15]), .Y(n131) );
  INVX2 U149 ( .A(B[16]), .Y(n132) );
  INVX2 U150 ( .A(B[17]), .Y(n133) );
  INVX2 U151 ( .A(B[18]), .Y(n134) );
  INVX2 U152 ( .A(B[19]), .Y(n135) );
  INVX2 U153 ( .A(B[20]), .Y(n136) );
  INVX2 U154 ( .A(B[21]), .Y(n137) );
  INVX2 U155 ( .A(B[22]), .Y(n138) );
  INVX2 U156 ( .A(B[23]), .Y(n139) );
  INVX2 U157 ( .A(B[24]), .Y(n140) );
  INVX2 U158 ( .A(B[25]), .Y(n141) );
  INVX2 U159 ( .A(B[26]), .Y(n142) );
  INVX2 U160 ( .A(B[27]), .Y(n143) );
  INVX2 U161 ( .A(B[28]), .Y(n144) );
  INVX2 U162 ( .A(B[29]), .Y(n145) );
  INVX2 U163 ( .A(B[30]), .Y(n146) );
  INVX2 U164 ( .A(B[9]), .Y(n147) );
  INVX2 U165 ( .A(B[10]), .Y(n148) );
  INVX2 U166 ( .A(A[2]), .Y(n149) );
  INVX2 U167 ( .A(B[8]), .Y(n150) );
  INVX2 U168 ( .A(A[1]), .Y(n151) );
  INVX2 U169 ( .A(A[3]), .Y(n152) );
  INVX2 U170 ( .A(A[4]), .Y(n153) );
  INVX2 U431 ( .A(A[5]), .Y(n154) );
  INVX2 U432 ( .A(A[6]), .Y(n155) );
endmodule


module CannyEdge_DW02_mult_21 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n17), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n18), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n16), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n22), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n21), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n34), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n35), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n37), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n38), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n39), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n33), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n34), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n35), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n36), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n37), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n38), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n39), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n33), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW01_cmp2_5 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180;

  MUX2X1 U60 ( .B(n60), .A(n61), .S(B[31]), .Y(LT_LE) );
  MUX2X1 U61 ( .B(n158), .A(n62), .S(A[31]), .Y(n61) );
  NAND2X1 U62 ( .A(A[30]), .B(n63), .Y(n62) );
  MUX2X1 U63 ( .B(n122), .A(TC), .S(A[31]), .Y(n60) );
  OAI21X1 U64 ( .A(B[31]), .B(n178), .C(n64), .Y(n63) );
  AOI21X1 U65 ( .A(A[29]), .B(n137), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n177), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n138), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n176), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n139), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n175), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n140), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n174), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n141), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n173), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n142), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n172), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n143), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n171), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n144), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n170), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n145), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n169), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n146), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n168), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n147), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n167), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n148), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n166), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n149), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n165), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n150), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n164), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n151), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n163), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n152), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n162), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n153), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n161), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n154), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n160), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n155), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n159), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n156), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n180), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n156), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n180), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n157), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n179), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n126), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n136), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n125), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n135), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n124), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n134), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n123), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n133), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n129), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n130), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n128), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n132), .C(n120), .Y(n119) );
  AOI22X1 U121 ( .A(n121), .B(A[0]), .C(A[1]), .D(n127), .Y(n120) );
  AOI21X1 U122 ( .A(B[1]), .B(n131), .C(B[0]), .Y(n121) );
  INVX2 U1 ( .A(n63), .Y(n122) );
  INVX2 U2 ( .A(B[4]), .Y(n123) );
  INVX2 U3 ( .A(B[5]), .Y(n124) );
  INVX2 U4 ( .A(B[6]), .Y(n125) );
  INVX2 U5 ( .A(B[7]), .Y(n126) );
  INVX2 U6 ( .A(B[1]), .Y(n127) );
  INVX2 U7 ( .A(B[2]), .Y(n128) );
  INVX2 U8 ( .A(B[3]), .Y(n129) );
  INVX2 U9 ( .A(A[3]), .Y(n130) );
  INVX2 U10 ( .A(A[1]), .Y(n131) );
  INVX2 U11 ( .A(A[2]), .Y(n132) );
  INVX2 U12 ( .A(A[4]), .Y(n133) );
  INVX2 U13 ( .A(A[5]), .Y(n134) );
  INVX2 U14 ( .A(A[6]), .Y(n135) );
  INVX2 U15 ( .A(A[7]), .Y(n136) );
  INVX2 U16 ( .A(B[29]), .Y(n137) );
  INVX2 U17 ( .A(B[28]), .Y(n138) );
  INVX2 U18 ( .A(B[27]), .Y(n139) );
  INVX2 U19 ( .A(B[26]), .Y(n140) );
  INVX2 U20 ( .A(B[25]), .Y(n141) );
  INVX2 U21 ( .A(B[24]), .Y(n142) );
  INVX2 U22 ( .A(B[23]), .Y(n143) );
  INVX2 U23 ( .A(B[22]), .Y(n144) );
  INVX2 U24 ( .A(B[21]), .Y(n145) );
  INVX2 U25 ( .A(B[20]), .Y(n146) );
  INVX2 U26 ( .A(B[19]), .Y(n147) );
  INVX2 U27 ( .A(B[18]), .Y(n148) );
  INVX2 U28 ( .A(B[17]), .Y(n149) );
  INVX2 U29 ( .A(B[16]), .Y(n150) );
  INVX2 U30 ( .A(B[15]), .Y(n151) );
  INVX2 U31 ( .A(B[14]), .Y(n152) );
  INVX2 U32 ( .A(B[13]), .Y(n153) );
  INVX2 U33 ( .A(B[12]), .Y(n154) );
  INVX2 U34 ( .A(B[11]), .Y(n155) );
  INVX2 U35 ( .A(B[10]), .Y(n156) );
  INVX2 U36 ( .A(B[8]), .Y(n157) );
  INVX2 U37 ( .A(TC), .Y(n158) );
  INVX2 U38 ( .A(A[11]), .Y(n159) );
  INVX2 U39 ( .A(A[12]), .Y(n160) );
  INVX2 U40 ( .A(A[13]), .Y(n161) );
  INVX2 U41 ( .A(A[14]), .Y(n162) );
  INVX2 U42 ( .A(A[15]), .Y(n163) );
  INVX2 U43 ( .A(A[16]), .Y(n164) );
  INVX2 U44 ( .A(A[17]), .Y(n165) );
  INVX2 U45 ( .A(A[18]), .Y(n166) );
  INVX2 U46 ( .A(A[19]), .Y(n167) );
  INVX2 U47 ( .A(A[20]), .Y(n168) );
  INVX2 U48 ( .A(A[21]), .Y(n169) );
  INVX2 U49 ( .A(A[22]), .Y(n170) );
  INVX2 U50 ( .A(A[23]), .Y(n171) );
  INVX2 U51 ( .A(A[24]), .Y(n172) );
  INVX2 U52 ( .A(A[25]), .Y(n173) );
  INVX2 U53 ( .A(A[26]), .Y(n174) );
  INVX2 U54 ( .A(A[27]), .Y(n175) );
  INVX2 U55 ( .A(A[28]), .Y(n176) );
  INVX2 U56 ( .A(A[29]), .Y(n177) );
  INVX2 U57 ( .A(A[30]), .Y(n178) );
  INVX2 U58 ( .A(A[8]), .Y(n179) );
  INVX2 U59 ( .A(A[9]), .Y(n180) );
endmodule


module CannyEdge_DW01_add_45 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_22 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \SUMB[7][7] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] ,
         \SUMB[5][1] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] ,
         \SUMB[4][1] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n60, n61, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign PRODUCT[1] = \ab[0][1] ;
  assign QA = TC;

  AND2X2 U2 ( .A(n41), .B(n66), .Y(n3) );
  AND2X2 U3 ( .A(n19), .B(n66), .Y(n4) );
  AND2X2 U4 ( .A(\ab[2][6] ), .B(n66), .Y(n5) );
  AND2X2 U5 ( .A(n28), .B(\SUMB[4][5] ), .Y(n6) );
  AND2X2 U6 ( .A(n26), .B(\SUMB[4][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[5][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n33), .B(\SUMB[2][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n34), .B(\SUMB[2][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n35), .B(\SUMB[2][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n36), .B(\SUMB[2][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n40), .B(\SUMB[6][1] ), .Y(n13) );
  AND2X2 U13 ( .A(n30), .B(\SUMB[6][2] ), .Y(n14) );
  AND2X2 U14 ( .A(n25), .B(\SUMB[6][4] ), .Y(n15) );
  AND2X2 U15 ( .A(n31), .B(\SUMB[6][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\SUMB[3][1] ), .B(n39), .Y(n17) );
  AND2X2 U17 ( .A(QA), .B(QB), .Y(n18) );
  AND2X2 U18 ( .A(n3), .B(n66), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[2][0] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][5] ), .B(\ab[0][7] ), .Y(n21) );
  AND2X2 U21 ( .A(n8), .B(\SUMB[6][3] ), .Y(n22) );
  AND2X2 U22 ( .A(n11), .B(\SUMB[3][4] ), .Y(n23) );
  AND2X2 U23 ( .A(n23), .B(\SUMB[4][4] ), .Y(n24) );
  AND2X2 U24 ( .A(n24), .B(\SUMB[5][4] ), .Y(n25) );
  AND2X2 U25 ( .A(n9), .B(\SUMB[3][2] ), .Y(n26) );
  AND2X2 U26 ( .A(n10), .B(\SUMB[3][3] ), .Y(n27) );
  AND2X2 U27 ( .A(n12), .B(\SUMB[3][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n27), .B(\SUMB[4][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n7), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n6), .B(\SUMB[5][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n21), .B(\SUMB[2][6] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[2][1] ), .B(\ab[0][3] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[2][2] ), .B(\ab[0][4] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[2][3] ), .B(\ab[0][5] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[2][4] ), .B(\ab[0][6] ), .Y(n36) );
  AND2X2 U36 ( .A(\SUMB[7][1] ), .B(n13), .Y(n37) );
  AND2X2 U37 ( .A(\SUMB[4][1] ), .B(n17), .Y(n38) );
  AND2X2 U38 ( .A(\SUMB[2][1] ), .B(n20), .Y(n39) );
  AND2X2 U39 ( .A(\SUMB[5][1] ), .B(n38), .Y(n40) );
  AND2X2 U40 ( .A(n32), .B(n5), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n66), .Y(n42) );
  AND2X2 U42 ( .A(n66), .B(n4), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n22), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n14), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n15), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n16), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n13), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n14), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n22), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n15), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n16), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n66), .B(n4), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n18), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\SUMB[7][0] ), .B(n66), .Y(\A1[5] ) );
  XOR2X1 U55 ( .A(\SUMB[2][1] ), .B(n20), .Y(\A1[1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][2] ), .B(n33), .Y(\SUMB[3][1] ) );
  XOR2X1 U57 ( .A(\SUMB[2][3] ), .B(n34), .Y(\SUMB[3][2] ) );
  XOR2X1 U58 ( .A(\SUMB[2][4] ), .B(n35), .Y(\SUMB[3][3] ) );
  XOR2X1 U59 ( .A(\SUMB[2][5] ), .B(n36), .Y(\SUMB[3][4] ) );
  XOR2X1 U60 ( .A(\SUMB[2][6] ), .B(n21), .Y(\SUMB[3][5] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n39), .Y(\A1[2] ) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n9), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n10), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n11), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n12), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(n5), .B(n32), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n17), .Y(\A1[3] ) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n26), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n27), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n23), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n28), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n66), .B(n41), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n38), .Y(\A1[4] ) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n7), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n29), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n24), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n6), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(n66), .B(n3), .Y(\SUMB[6][5] ) );
  XOR2X1 U79 ( .A(\SUMB[6][1] ), .B(n40), .Y(\SUMB[7][0] ) );
  XOR2X1 U80 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U81 ( .A(\SUMB[6][3] ), .B(n8), .Y(\SUMB[7][2] ) );
  XOR2X1 U82 ( .A(\SUMB[6][4] ), .B(n25), .Y(\SUMB[7][3] ) );
  XOR2X1 U83 ( .A(\SUMB[6][5] ), .B(n31), .Y(\SUMB[7][4] ) );
  XOR2X1 U84 ( .A(n66), .B(n19), .Y(\SUMB[7][5] ) );
  XOR2X1 U85 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  XOR2X1 U86 ( .A(\ab[0][2] ), .B(\ab[2][0] ), .Y(\A1[0] ) );
  XOR2X1 U87 ( .A(\ab[0][3] ), .B(\ab[2][1] ), .Y(\SUMB[2][1] ) );
  XOR2X1 U88 ( .A(\ab[0][4] ), .B(\ab[2][2] ), .Y(\SUMB[2][2] ) );
  XOR2X1 U89 ( .A(\ab[0][5] ), .B(\ab[2][3] ), .Y(\SUMB[2][3] ) );
  XOR2X1 U90 ( .A(\ab[0][6] ), .B(\ab[2][4] ), .Y(\SUMB[2][4] ) );
  XOR2X1 U91 ( .A(\ab[0][7] ), .B(\ab[2][5] ), .Y(\SUMB[2][5] ) );
  XOR2X1 U92 ( .A(n66), .B(\ab[2][6] ), .Y(\SUMB[2][6] ) );
  NOR2X1 U104 ( .A(n65), .B(n72), .Y(\ab[2][6] ) );
  NOR2X1 U105 ( .A(n65), .B(n71), .Y(\ab[2][5] ) );
  NOR2X1 U106 ( .A(n65), .B(n70), .Y(\ab[2][4] ) );
  NOR2X1 U107 ( .A(n65), .B(n69), .Y(\ab[2][3] ) );
  NOR2X1 U108 ( .A(n65), .B(n68), .Y(\ab[2][2] ) );
  NOR2X1 U109 ( .A(n65), .B(n67), .Y(\ab[2][1] ) );
  NOR2X1 U110 ( .A(n65), .B(n74), .Y(\ab[2][0] ) );
  MUX2X1 U111 ( .B(n60), .A(n61), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U112 ( .A(B[7]), .B(n65), .Y(n61) );
  NOR2X1 U113 ( .A(n72), .B(n73), .Y(\ab[0][6] ) );
  NOR2X1 U114 ( .A(n71), .B(n73), .Y(\ab[0][5] ) );
  NOR2X1 U115 ( .A(n70), .B(n73), .Y(\ab[0][4] ) );
  NOR2X1 U116 ( .A(n69), .B(n73), .Y(\ab[0][3] ) );
  NOR2X1 U117 ( .A(n68), .B(n73), .Y(\ab[0][2] ) );
  NOR2X1 U118 ( .A(n67), .B(n73), .Y(\ab[0][1] ) );
  NAND2X1 U119 ( .A(QA), .B(B[7]), .Y(n60) );
  NOR2X1 U120 ( .A(B[7]), .B(n65), .Y(QB) );
  NOR2X1 U121 ( .A(n74), .B(n73), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_45 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n37, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n65) );
  INVX2 U97 ( .A(n60), .Y(n66) );
  INVX2 U98 ( .A(B[1]), .Y(n67) );
  INVX2 U99 ( .A(B[2]), .Y(n68) );
  INVX2 U100 ( .A(B[3]), .Y(n69) );
  INVX2 U101 ( .A(B[4]), .Y(n70) );
  INVX2 U102 ( .A(B[5]), .Y(n71) );
  INVX2 U103 ( .A(B[6]), .Y(n72) );
  INVX2 U122 ( .A(A[0]), .Y(n73) );
  INVX2 U123 ( .A(B[0]), .Y(n74) );
endmodule


module CannyEdge_DW01_add_47 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_23 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] ,
         \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] ,
         \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] ,
         \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n57, n58, n61, n62;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign PRODUCT[0] = \ab[2][0] ;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n23), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n22), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n21), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n20), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n19), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n18), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n24), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(\SUMB[7][7] ), .B(n5), .Y(n3) );
  AND2X2 U3 ( .A(n28), .B(n62), .Y(n4) );
  AND2X2 U4 ( .A(n27), .B(n62), .Y(n5) );
  AND2X2 U5 ( .A(n44), .B(\SUMB[3][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n45), .B(\SUMB[3][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n46), .B(\SUMB[3][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n47), .B(\SUMB[3][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n43), .B(\SUMB[3][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n42), .B(\SUMB[6][1] ), .Y(n11) );
  AND2X2 U11 ( .A(n34), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n35), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n36), .B(\SUMB[6][4] ), .Y(n14) );
  AND2X2 U14 ( .A(n37), .B(\SUMB[6][5] ), .Y(n15) );
  AND2X2 U15 ( .A(n39), .B(\SUMB[6][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\SUMB[4][1] ), .B(n41), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][6] ), .B(\ab[1][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][5] ), .B(\ab[1][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][4] ), .B(\ab[1][3] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][3] ), .B(\ab[1][2] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][2] ), .B(\ab[1][1] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[2][1] ), .B(\ab[1][0] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[2][7] ), .B(\ab[1][6] ), .Y(n24) );
  AND2X2 U24 ( .A(QA), .B(QB), .Y(n25) );
  AND2X2 U25 ( .A(n4), .B(n62), .Y(n26) );
  AND2X2 U26 ( .A(n26), .B(n62), .Y(n27) );
  AND2X2 U27 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n28) );
  AND2X2 U28 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n29) );
  AND2X2 U29 ( .A(n6), .B(\SUMB[4][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n7), .B(\SUMB[4][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n8), .B(\SUMB[4][4] ), .Y(n32) );
  AND2X2 U32 ( .A(n9), .B(\SUMB[4][5] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][2] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][3] ), .Y(n35) );
  AND2X2 U35 ( .A(n32), .B(\SUMB[5][4] ), .Y(n36) );
  AND2X2 U36 ( .A(n33), .B(\SUMB[5][5] ), .Y(n37) );
  AND2X2 U37 ( .A(n10), .B(\SUMB[4][6] ), .Y(n38) );
  AND2X2 U38 ( .A(n38), .B(\SUMB[5][6] ), .Y(n39) );
  AND2X2 U39 ( .A(\SUMB[7][1] ), .B(n11), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[3][1] ), .B(n29), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[5][1] ), .B(n17), .Y(n42) );
  AND2X2 U42 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n43) );
  AND2X2 U43 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n44) );
  AND2X2 U44 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n45) );
  AND2X2 U45 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n46) );
  AND2X2 U46 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][0] ), .B(n62), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][6] ), .B(n16), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][3] ), .B(n13), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][5] ), .B(n15), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][2] ), .B(n12), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][4] ), .B(n14), .Y(n53) );
  XOR2X1 U53 ( .A(\SUMB[7][1] ), .B(n11), .Y(\A1[6] ) );
  XOR2X1 U54 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U55 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U56 ( .A(\SUMB[7][4] ), .B(n14), .Y(\A1[9] ) );
  XOR2X1 U57 ( .A(\SUMB[7][5] ), .B(n15), .Y(\A1[10] ) );
  XOR2X1 U58 ( .A(\SUMB[7][6] ), .B(n16), .Y(\A1[11] ) );
  XOR2X1 U59 ( .A(\SUMB[7][7] ), .B(n5), .Y(\A1[12] ) );
  XOR2X1 U60 ( .A(n25), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U61 ( .A(\ab[1][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U62 ( .A(\ab[1][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U63 ( .A(\ab[1][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U64 ( .A(\ab[1][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U65 ( .A(\ab[1][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U66 ( .A(\ab[1][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U67 ( .A(\ab[1][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U68 ( .A(\SUMB[7][0] ), .B(n62), .Y(\A1[5] ) );
  XOR2X1 U69 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U70 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U71 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U72 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U73 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U74 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U75 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U76 ( .A(\SUMB[3][1] ), .B(n29), .Y(\A1[2] ) );
  XOR2X1 U77 ( .A(\SUMB[3][2] ), .B(n44), .Y(\SUMB[4][1] ) );
  XOR2X1 U78 ( .A(\SUMB[3][3] ), .B(n45), .Y(\SUMB[4][2] ) );
  XOR2X1 U79 ( .A(\SUMB[3][4] ), .B(n46), .Y(\SUMB[4][3] ) );
  XOR2X1 U80 ( .A(\SUMB[3][5] ), .B(n47), .Y(\SUMB[4][4] ) );
  XOR2X1 U81 ( .A(\SUMB[3][6] ), .B(n43), .Y(\SUMB[4][5] ) );
  XOR2X1 U82 ( .A(n62), .B(n28), .Y(\SUMB[4][6] ) );
  XOR2X1 U83 ( .A(\SUMB[4][1] ), .B(n41), .Y(\A1[3] ) );
  XOR2X1 U84 ( .A(\SUMB[4][2] ), .B(n6), .Y(\SUMB[5][1] ) );
  XOR2X1 U85 ( .A(\SUMB[4][3] ), .B(n7), .Y(\SUMB[5][2] ) );
  XOR2X1 U86 ( .A(\SUMB[4][4] ), .B(n8), .Y(\SUMB[5][3] ) );
  XOR2X1 U87 ( .A(\SUMB[4][5] ), .B(n9), .Y(\SUMB[5][4] ) );
  XOR2X1 U88 ( .A(\SUMB[4][6] ), .B(n10), .Y(\SUMB[5][5] ) );
  XOR2X1 U89 ( .A(n62), .B(n4), .Y(\SUMB[5][6] ) );
  XOR2X1 U90 ( .A(\SUMB[5][1] ), .B(n17), .Y(\A1[4] ) );
  XOR2X1 U91 ( .A(\SUMB[5][2] ), .B(n30), .Y(\SUMB[6][1] ) );
  XOR2X1 U92 ( .A(\SUMB[5][3] ), .B(n31), .Y(\SUMB[6][2] ) );
  XOR2X1 U93 ( .A(\SUMB[5][4] ), .B(n32), .Y(\SUMB[6][3] ) );
  XOR2X1 U94 ( .A(\SUMB[5][5] ), .B(n33), .Y(\SUMB[6][4] ) );
  XOR2X1 U95 ( .A(\SUMB[5][6] ), .B(n38), .Y(\SUMB[6][5] ) );
  XOR2X1 U96 ( .A(n62), .B(n26), .Y(\SUMB[6][6] ) );
  XOR2X1 U97 ( .A(\SUMB[6][1] ), .B(n42), .Y(\SUMB[7][0] ) );
  XOR2X1 U98 ( .A(\SUMB[6][2] ), .B(n34), .Y(\SUMB[7][1] ) );
  XOR2X1 U99 ( .A(\SUMB[6][3] ), .B(n35), .Y(\SUMB[7][2] ) );
  XOR2X1 U100 ( .A(\SUMB[6][4] ), .B(n36), .Y(\SUMB[7][3] ) );
  XOR2X1 U101 ( .A(\SUMB[6][5] ), .B(n37), .Y(\SUMB[7][4] ) );
  XOR2X1 U102 ( .A(\SUMB[6][6] ), .B(n39), .Y(\SUMB[7][5] ) );
  XOR2X1 U103 ( .A(n62), .B(n27), .Y(\SUMB[7][6] ) );
  XOR2X1 U104 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  MUX2X1 U107 ( .B(n57), .A(n58), .S(A[1]), .Y(\ab[1][7] ) );
  AND2X1 U108 ( .A(B[6]), .B(A[1]), .Y(\ab[1][6] ) );
  AND2X1 U109 ( .A(B[5]), .B(A[1]), .Y(\ab[1][5] ) );
  AND2X1 U110 ( .A(B[4]), .B(A[1]), .Y(\ab[1][4] ) );
  AND2X1 U111 ( .A(B[3]), .B(A[1]), .Y(\ab[1][3] ) );
  AND2X1 U112 ( .A(B[2]), .B(A[1]), .Y(\ab[1][2] ) );
  AND2X1 U113 ( .A(B[1]), .B(A[1]), .Y(\ab[1][1] ) );
  AND2X1 U114 ( .A(B[0]), .B(A[1]), .Y(\ab[1][0] ) );
  MUX2X1 U115 ( .B(n57), .A(n58), .S(A[2]), .Y(\ab[2][7] ) );
  NAND2X1 U116 ( .A(B[7]), .B(n61), .Y(n58) );
  AND2X1 U117 ( .A(B[6]), .B(A[2]), .Y(\ab[2][6] ) );
  AND2X1 U118 ( .A(B[5]), .B(A[2]), .Y(\ab[2][5] ) );
  AND2X1 U119 ( .A(B[4]), .B(A[2]), .Y(\ab[2][4] ) );
  AND2X1 U120 ( .A(B[3]), .B(A[2]), .Y(\ab[2][3] ) );
  AND2X1 U121 ( .A(B[2]), .B(A[2]), .Y(\ab[2][2] ) );
  AND2X1 U122 ( .A(B[1]), .B(A[2]), .Y(\ab[2][1] ) );
  NAND2X1 U123 ( .A(QA), .B(B[7]), .Y(n57) );
  NOR2X1 U124 ( .A(B[7]), .B(n61), .Y(QB) );
  AND2X1 U125 ( .A(B[0]), .B(A[2]), .Y(\ab[2][0] ) );
  CannyEdge_DW01_add_47 FS_1 ( .A({\A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({n3, n49, n51, n53, n50, n52, n40, n48, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U126 ( .A(QA), .Y(n61) );
  INVX2 U127 ( .A(n57), .Y(n62) );
endmodule


module CannyEdge_DW01_cmp2_6 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188;

  MUX2X1 U63 ( .B(n63), .A(n64), .S(B[31]), .Y(LT_LE) );
  MUX2X1 U64 ( .B(n160), .A(n65), .S(A[31]), .Y(n64) );
  NOR2X1 U65 ( .A(n66), .B(n186), .Y(n65) );
  MUX2X1 U66 ( .B(n67), .A(TC), .S(A[31]), .Y(n63) );
  NAND2X1 U67 ( .A(n66), .B(n186), .Y(n67) );
  AOI21X1 U68 ( .A(n134), .B(B[29]), .C(n127), .Y(n66) );
  OAI21X1 U69 ( .A(B[29]), .B(n134), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(A[28]), .B(n185), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(B[28]), .B(n135), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(A[27]), .B(n184), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(B[27]), .B(n136), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(A[26]), .B(n183), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(B[26]), .B(n137), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(A[25]), .B(n182), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(B[25]), .B(n138), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(A[24]), .B(n181), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(B[24]), .B(n139), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(A[23]), .B(n180), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(B[23]), .B(n140), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(A[22]), .B(n179), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(B[22]), .B(n141), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(A[21]), .B(n178), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(B[21]), .B(n142), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(A[20]), .B(n177), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(B[20]), .B(n143), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(A[19]), .B(n176), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(B[19]), .B(n144), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(A[18]), .B(n175), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(B[18]), .B(n145), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(A[17]), .B(n174), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(B[17]), .B(n146), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(A[16]), .B(n173), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(B[16]), .B(n147), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(A[15]), .B(n172), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(B[15]), .B(n148), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(A[14]), .B(n171), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(B[14]), .B(n149), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(A[13]), .B(n170), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(B[13]), .B(n150), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(A[12]), .B(n169), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(B[12]), .B(n151), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(A[11]), .B(n168), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(B[11]), .B(n152), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(A[10]), .B(n167), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(B[10]), .B(n153), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(A[9]), .B(n188), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(B[9]), .B(n154), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(A[8]), .B(n187), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(B[8]), .B(n155), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(A[7]), .B(n161), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(B[7]), .B(n156), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(A[6]), .B(n162), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(B[6]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(A[5]), .B(n163), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(B[5]), .B(n158), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(A[4]), .B(n164), .C(n118), .Y(n117) );
  AOI21X1 U119 ( .A(B[4]), .B(n159), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(A[3]), .B(n133), .C(n120), .Y(n119) );
  OAI21X1 U121 ( .A(B[3]), .B(n131), .C(n121), .Y(n120) );
  AOI21X1 U122 ( .A(A[2]), .B(n165), .C(n122), .Y(n121) );
  AOI21X1 U123 ( .A(B[2]), .B(n130), .C(n123), .Y(n122) );
  OAI21X1 U124 ( .A(A[1]), .B(n132), .C(n124), .Y(n123) );
  OAI21X1 U125 ( .A(B[1]), .B(n129), .C(n125), .Y(n124) );
  AOI21X1 U126 ( .A(A[0]), .B(n166), .C(n126), .Y(n125) );
  AOI21X1 U127 ( .A(B[0]), .B(n128), .C(LEQ), .Y(n126) );
  INVX2 U1 ( .A(n68), .Y(n127) );
  INVX2 U2 ( .A(A[0]), .Y(n128) );
  INVX2 U3 ( .A(A[1]), .Y(n129) );
  INVX2 U4 ( .A(A[2]), .Y(n130) );
  INVX2 U5 ( .A(A[3]), .Y(n131) );
  INVX2 U6 ( .A(B[1]), .Y(n132) );
  INVX2 U7 ( .A(B[3]), .Y(n133) );
  INVX2 U8 ( .A(A[29]), .Y(n134) );
  INVX2 U9 ( .A(A[28]), .Y(n135) );
  INVX2 U10 ( .A(A[27]), .Y(n136) );
  INVX2 U11 ( .A(A[26]), .Y(n137) );
  INVX2 U12 ( .A(A[25]), .Y(n138) );
  INVX2 U13 ( .A(A[24]), .Y(n139) );
  INVX2 U14 ( .A(A[23]), .Y(n140) );
  INVX2 U15 ( .A(A[22]), .Y(n141) );
  INVX2 U16 ( .A(A[21]), .Y(n142) );
  INVX2 U17 ( .A(A[20]), .Y(n143) );
  INVX2 U18 ( .A(A[19]), .Y(n144) );
  INVX2 U19 ( .A(A[18]), .Y(n145) );
  INVX2 U20 ( .A(A[17]), .Y(n146) );
  INVX2 U21 ( .A(A[16]), .Y(n147) );
  INVX2 U22 ( .A(A[15]), .Y(n148) );
  INVX2 U23 ( .A(A[14]), .Y(n149) );
  INVX2 U24 ( .A(A[13]), .Y(n150) );
  INVX2 U25 ( .A(A[12]), .Y(n151) );
  INVX2 U26 ( .A(A[11]), .Y(n152) );
  INVX2 U27 ( .A(A[10]), .Y(n153) );
  INVX2 U28 ( .A(A[9]), .Y(n154) );
  INVX2 U29 ( .A(A[8]), .Y(n155) );
  INVX2 U30 ( .A(A[7]), .Y(n156) );
  INVX2 U31 ( .A(A[6]), .Y(n157) );
  INVX2 U32 ( .A(A[5]), .Y(n158) );
  INVX2 U33 ( .A(A[4]), .Y(n159) );
  INVX2 U34 ( .A(TC), .Y(n160) );
  INVX2 U35 ( .A(B[7]), .Y(n161) );
  INVX2 U36 ( .A(B[6]), .Y(n162) );
  INVX2 U37 ( .A(B[5]), .Y(n163) );
  INVX2 U38 ( .A(B[4]), .Y(n164) );
  INVX2 U39 ( .A(B[2]), .Y(n165) );
  INVX2 U40 ( .A(B[0]), .Y(n166) );
  INVX2 U41 ( .A(B[10]), .Y(n167) );
  INVX2 U42 ( .A(B[11]), .Y(n168) );
  INVX2 U43 ( .A(B[12]), .Y(n169) );
  INVX2 U44 ( .A(B[13]), .Y(n170) );
  INVX2 U45 ( .A(B[14]), .Y(n171) );
  INVX2 U46 ( .A(B[15]), .Y(n172) );
  INVX2 U47 ( .A(B[16]), .Y(n173) );
  INVX2 U48 ( .A(B[17]), .Y(n174) );
  INVX2 U49 ( .A(B[18]), .Y(n175) );
  INVX2 U50 ( .A(B[19]), .Y(n176) );
  INVX2 U51 ( .A(B[20]), .Y(n177) );
  INVX2 U52 ( .A(B[21]), .Y(n178) );
  INVX2 U53 ( .A(B[22]), .Y(n179) );
  INVX2 U54 ( .A(B[23]), .Y(n180) );
  INVX2 U55 ( .A(B[24]), .Y(n181) );
  INVX2 U56 ( .A(B[25]), .Y(n182) );
  INVX2 U57 ( .A(B[26]), .Y(n183) );
  INVX2 U58 ( .A(B[27]), .Y(n184) );
  INVX2 U59 ( .A(B[28]), .Y(n185) );
  INVX2 U60 ( .A(B[30]), .Y(n186) );
  INVX2 U61 ( .A(B[8]), .Y(n187) );
  INVX2 U62 ( .A(B[9]), .Y(n188) );
endmodule


module CannyEdge_DW01_addsub_16 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  AND2X2 U1 ( .A(n12), .B(B_AS[29]), .Y(n1) );
  AND2X2 U2 ( .A(n13), .B(B_AS[27]), .Y(n2) );
  AND2X2 U3 ( .A(n14), .B(B_AS[25]), .Y(n3) );
  AND2X2 U4 ( .A(n15), .B(B_AS[23]), .Y(n4) );
  AND2X2 U5 ( .A(n16), .B(B_AS[21]), .Y(n5) );
  AND2X2 U6 ( .A(n17), .B(B_AS[19]), .Y(n6) );
  AND2X2 U7 ( .A(n18), .B(B_AS[17]), .Y(n7) );
  AND2X2 U8 ( .A(n19), .B(B_AS[15]), .Y(n8) );
  AND2X2 U9 ( .A(n20), .B(B_AS[13]), .Y(n9) );
  AND2X2 U10 ( .A(n21), .B(B_AS[11]), .Y(n10) );
  AND2X2 U11 ( .A(n22), .B(B_AS[9]), .Y(n11) );
  AND2X2 U12 ( .A(n2), .B(B_AS[28]), .Y(n12) );
  AND2X2 U13 ( .A(n3), .B(B_AS[26]), .Y(n13) );
  AND2X2 U14 ( .A(n4), .B(B_AS[24]), .Y(n14) );
  AND2X2 U15 ( .A(n5), .B(B_AS[22]), .Y(n15) );
  AND2X2 U16 ( .A(n6), .B(B_AS[20]), .Y(n16) );
  AND2X2 U17 ( .A(n7), .B(B_AS[18]), .Y(n17) );
  AND2X2 U18 ( .A(n8), .B(B_AS[16]), .Y(n18) );
  AND2X2 U19 ( .A(n9), .B(B_AS[14]), .Y(n19) );
  AND2X2 U20 ( .A(n10), .B(B_AS[12]), .Y(n20) );
  AND2X2 U21 ( .A(n11), .B(B_AS[10]), .Y(n21) );
  AND2X2 U22 ( .A(carry[8]), .B(B_AS[8]), .Y(n22) );
  AND2X2 U23 ( .A(n1), .B(B_AS[30]), .Y(n23) );
  XOR2X1 U24 ( .A(B_AS[31]), .B(n23), .Y(SUM[31]) );
  XOR2X1 U25 ( .A(n1), .B(B_AS[30]), .Y(SUM[30]) );
  XOR2X1 U26 ( .A(n12), .B(B_AS[29]), .Y(SUM[29]) );
  XOR2X1 U27 ( .A(n2), .B(B_AS[28]), .Y(SUM[28]) );
  XOR2X1 U28 ( .A(n13), .B(B_AS[27]), .Y(SUM[27]) );
  XOR2X1 U29 ( .A(n3), .B(B_AS[26]), .Y(SUM[26]) );
  XOR2X1 U30 ( .A(n14), .B(B_AS[25]), .Y(SUM[25]) );
  XOR2X1 U31 ( .A(n4), .B(B_AS[24]), .Y(SUM[24]) );
  XOR2X1 U32 ( .A(n15), .B(B_AS[23]), .Y(SUM[23]) );
  XOR2X1 U33 ( .A(n5), .B(B_AS[22]), .Y(SUM[22]) );
  XOR2X1 U34 ( .A(n16), .B(B_AS[21]), .Y(SUM[21]) );
  XOR2X1 U35 ( .A(n6), .B(B_AS[20]), .Y(SUM[20]) );
  XOR2X1 U36 ( .A(n17), .B(B_AS[19]), .Y(SUM[19]) );
  XOR2X1 U37 ( .A(n7), .B(B_AS[18]), .Y(SUM[18]) );
  XOR2X1 U38 ( .A(n18), .B(B_AS[17]), .Y(SUM[17]) );
  XOR2X1 U39 ( .A(n8), .B(B_AS[16]), .Y(SUM[16]) );
  XOR2X1 U40 ( .A(n19), .B(B_AS[15]), .Y(SUM[15]) );
  XOR2X1 U41 ( .A(n9), .B(B_AS[14]), .Y(SUM[14]) );
  XOR2X1 U42 ( .A(n20), .B(B_AS[13]), .Y(SUM[13]) );
  XOR2X1 U43 ( .A(n10), .B(B_AS[12]), .Y(SUM[12]) );
  XOR2X1 U44 ( .A(n21), .B(B_AS[11]), .Y(SUM[11]) );
  XOR2X1 U45 ( .A(n11), .B(B_AS[10]), .Y(SUM[10]) );
  XOR2X1 U46 ( .A(n22), .B(B_AS[9]), .Y(SUM[9]) );
  XOR2X1 U47 ( .A(carry[8]), .B(B_AS[8]), .Y(SUM[8]) );
  XOR2X1 U48 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U49 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U50 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U51 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U52 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U53 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U54 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U55 ( .A(B[31]), .B(carry[0]), .Y(B_AS[31]) );
  XOR2X1 U56 ( .A(B[30]), .B(carry[0]), .Y(B_AS[30]) );
  XOR2X1 U57 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U58 ( .A(B[29]), .B(carry[0]), .Y(B_AS[29]) );
  XOR2X1 U59 ( .A(B[28]), .B(carry[0]), .Y(B_AS[28]) );
  XOR2X1 U60 ( .A(B[27]), .B(carry[0]), .Y(B_AS[27]) );
  XOR2X1 U61 ( .A(B[26]), .B(carry[0]), .Y(B_AS[26]) );
  XOR2X1 U62 ( .A(B[25]), .B(carry[0]), .Y(B_AS[25]) );
  XOR2X1 U63 ( .A(B[24]), .B(carry[0]), .Y(B_AS[24]) );
  XOR2X1 U64 ( .A(B[23]), .B(carry[0]), .Y(B_AS[23]) );
  XOR2X1 U65 ( .A(B[22]), .B(carry[0]), .Y(B_AS[22]) );
  XOR2X1 U66 ( .A(B[21]), .B(carry[0]), .Y(B_AS[21]) );
  XOR2X1 U67 ( .A(B[20]), .B(carry[0]), .Y(B_AS[20]) );
  XOR2X1 U68 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U69 ( .A(B[19]), .B(carry[0]), .Y(B_AS[19]) );
  XOR2X1 U70 ( .A(B[18]), .B(carry[0]), .Y(B_AS[18]) );
  XOR2X1 U71 ( .A(B[17]), .B(carry[0]), .Y(B_AS[17]) );
  XOR2X1 U72 ( .A(B[16]), .B(carry[0]), .Y(B_AS[16]) );
  XOR2X1 U73 ( .A(B[15]), .B(carry[0]), .Y(B_AS[15]) );
  XOR2X1 U74 ( .A(B[14]), .B(carry[0]), .Y(B_AS[14]) );
  XOR2X1 U75 ( .A(B[13]), .B(carry[0]), .Y(B_AS[13]) );
  XOR2X1 U76 ( .A(B[12]), .B(carry[0]), .Y(B_AS[12]) );
  XOR2X1 U77 ( .A(B[11]), .B(carry[0]), .Y(B_AS[11]) );
  XOR2X1 U78 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U79 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_add_48 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140;
  assign SUM[6] = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2X1 U2 ( .A(n126), .B(B[7]), .Y(SUM[7]) );
  NAND2X1 U29 ( .A(A[7]), .B(B[7]), .Y(n114) );
  XOR2X1 U30 ( .A(n28), .B(n29), .Y(SUM[9]) );
  NOR2X1 U31 ( .A(n122), .B(n30), .Y(n29) );
  XOR2X1 U32 ( .A(n32), .B(n114), .Y(SUM[8]) );
  NAND2X1 U33 ( .A(n125), .B(n33), .Y(n32) );
  XOR2X1 U34 ( .A(n35), .B(n36), .Y(SUM[29]) );
  XOR2X1 U35 ( .A(B[29]), .B(A[29]), .Y(n36) );
  OAI21X1 U36 ( .A(n37), .B(n38), .C(n39), .Y(n35) );
  XOR2X1 U37 ( .A(n40), .B(n38), .Y(SUM[28]) );
  AOI21X1 U38 ( .A(n128), .B(n41), .C(n42), .Y(n38) );
  NAND2X1 U39 ( .A(n127), .B(n39), .Y(n40) );
  NAND2X1 U40 ( .A(B[28]), .B(A[28]), .Y(n39) );
  NOR2X1 U41 ( .A(B[28]), .B(A[28]), .Y(n37) );
  XOR2X1 U42 ( .A(n41), .B(n44), .Y(SUM[27]) );
  NOR2X1 U43 ( .A(n42), .B(n43), .Y(n44) );
  NOR2X1 U44 ( .A(B[27]), .B(A[27]), .Y(n43) );
  AND2X1 U45 ( .A(B[27]), .B(A[27]), .Y(n42) );
  OAI21X1 U46 ( .A(n45), .B(n46), .C(n47), .Y(n41) );
  XOR2X1 U47 ( .A(n48), .B(n46), .Y(SUM[26]) );
  AOI21X1 U48 ( .A(n130), .B(n49), .C(n50), .Y(n46) );
  NAND2X1 U49 ( .A(n129), .B(n47), .Y(n48) );
  NAND2X1 U50 ( .A(B[26]), .B(A[26]), .Y(n47) );
  NOR2X1 U51 ( .A(B[26]), .B(A[26]), .Y(n45) );
  XOR2X1 U52 ( .A(n49), .B(n52), .Y(SUM[25]) );
  NOR2X1 U53 ( .A(n50), .B(n51), .Y(n52) );
  NOR2X1 U54 ( .A(B[25]), .B(A[25]), .Y(n51) );
  AND2X1 U55 ( .A(B[25]), .B(A[25]), .Y(n50) );
  OAI21X1 U56 ( .A(n53), .B(n54), .C(n55), .Y(n49) );
  XOR2X1 U57 ( .A(n56), .B(n54), .Y(SUM[24]) );
  AOI21X1 U58 ( .A(n132), .B(n57), .C(n58), .Y(n54) );
  NAND2X1 U59 ( .A(n131), .B(n55), .Y(n56) );
  NAND2X1 U60 ( .A(B[24]), .B(A[24]), .Y(n55) );
  NOR2X1 U61 ( .A(B[24]), .B(A[24]), .Y(n53) );
  XOR2X1 U62 ( .A(n57), .B(n60), .Y(SUM[23]) );
  NOR2X1 U63 ( .A(n58), .B(n59), .Y(n60) );
  NOR2X1 U64 ( .A(B[23]), .B(A[23]), .Y(n59) );
  AND2X1 U65 ( .A(B[23]), .B(A[23]), .Y(n58) );
  OAI21X1 U66 ( .A(n61), .B(n62), .C(n63), .Y(n57) );
  XOR2X1 U67 ( .A(n64), .B(n62), .Y(SUM[22]) );
  AOI21X1 U68 ( .A(n134), .B(n65), .C(n66), .Y(n62) );
  NAND2X1 U69 ( .A(n133), .B(n63), .Y(n64) );
  NAND2X1 U70 ( .A(B[22]), .B(A[22]), .Y(n63) );
  NOR2X1 U71 ( .A(B[22]), .B(A[22]), .Y(n61) );
  XOR2X1 U72 ( .A(n65), .B(n68), .Y(SUM[21]) );
  NOR2X1 U73 ( .A(n66), .B(n67), .Y(n68) );
  NOR2X1 U74 ( .A(B[21]), .B(A[21]), .Y(n67) );
  AND2X1 U75 ( .A(B[21]), .B(A[21]), .Y(n66) );
  OAI21X1 U76 ( .A(n69), .B(n70), .C(n71), .Y(n65) );
  XOR2X1 U77 ( .A(n72), .B(n70), .Y(SUM[20]) );
  AOI21X1 U78 ( .A(n136), .B(n73), .C(n74), .Y(n70) );
  NAND2X1 U79 ( .A(n135), .B(n71), .Y(n72) );
  NAND2X1 U80 ( .A(B[20]), .B(A[20]), .Y(n71) );
  NOR2X1 U81 ( .A(B[20]), .B(A[20]), .Y(n69) );
  XOR2X1 U82 ( .A(n73), .B(n76), .Y(SUM[19]) );
  NOR2X1 U83 ( .A(n74), .B(n75), .Y(n76) );
  NOR2X1 U84 ( .A(B[19]), .B(A[19]), .Y(n75) );
  AND2X1 U85 ( .A(B[19]), .B(A[19]), .Y(n74) );
  OAI21X1 U86 ( .A(n77), .B(n78), .C(n79), .Y(n73) );
  XOR2X1 U87 ( .A(n80), .B(n78), .Y(SUM[18]) );
  AOI21X1 U88 ( .A(n138), .B(n81), .C(n82), .Y(n78) );
  NAND2X1 U89 ( .A(n137), .B(n79), .Y(n80) );
  NAND2X1 U90 ( .A(B[18]), .B(A[18]), .Y(n79) );
  NOR2X1 U91 ( .A(B[18]), .B(A[18]), .Y(n77) );
  XOR2X1 U92 ( .A(n81), .B(n84), .Y(SUM[17]) );
  NOR2X1 U93 ( .A(n82), .B(n83), .Y(n84) );
  NOR2X1 U94 ( .A(B[17]), .B(A[17]), .Y(n83) );
  AND2X1 U95 ( .A(B[17]), .B(A[17]), .Y(n82) );
  OAI21X1 U96 ( .A(n85), .B(n86), .C(n87), .Y(n81) );
  XOR2X1 U97 ( .A(n88), .B(n86), .Y(SUM[16]) );
  AOI21X1 U98 ( .A(n140), .B(n89), .C(n90), .Y(n86) );
  NAND2X1 U99 ( .A(n139), .B(n87), .Y(n88) );
  NAND2X1 U100 ( .A(B[16]), .B(A[16]), .Y(n87) );
  NOR2X1 U101 ( .A(B[16]), .B(A[16]), .Y(n85) );
  XOR2X1 U102 ( .A(n89), .B(n92), .Y(SUM[15]) );
  NOR2X1 U103 ( .A(n90), .B(n91), .Y(n92) );
  NOR2X1 U104 ( .A(B[15]), .B(A[15]), .Y(n91) );
  AND2X1 U105 ( .A(B[15]), .B(A[15]), .Y(n90) );
  OAI21X1 U106 ( .A(n93), .B(n94), .C(n95), .Y(n89) );
  XOR2X1 U107 ( .A(n96), .B(n94), .Y(SUM[14]) );
  AOI21X1 U108 ( .A(n116), .B(n97), .C(n98), .Y(n94) );
  NAND2X1 U109 ( .A(n115), .B(n95), .Y(n96) );
  NAND2X1 U110 ( .A(B[14]), .B(A[14]), .Y(n95) );
  NOR2X1 U111 ( .A(B[14]), .B(A[14]), .Y(n93) );
  XOR2X1 U112 ( .A(n97), .B(n100), .Y(SUM[13]) );
  NOR2X1 U113 ( .A(n98), .B(n99), .Y(n100) );
  NOR2X1 U114 ( .A(B[13]), .B(A[13]), .Y(n99) );
  AND2X1 U115 ( .A(B[13]), .B(A[13]), .Y(n98) );
  OAI21X1 U116 ( .A(n101), .B(n118), .C(n102), .Y(n97) );
  XOR2X1 U117 ( .A(n103), .B(n118), .Y(SUM[12]) );
  OAI21X1 U118 ( .A(n105), .B(n106), .C(n107), .Y(n104) );
  AOI21X1 U119 ( .A(n108), .B(n121), .C(n120), .Y(n106) );
  NAND2X1 U120 ( .A(n117), .B(n102), .Y(n103) );
  NAND2X1 U121 ( .A(B[12]), .B(A[12]), .Y(n102) );
  NOR2X1 U122 ( .A(B[12]), .B(A[12]), .Y(n101) );
  XOR2X1 U123 ( .A(n110), .B(n111), .Y(SUM[11]) );
  NOR2X1 U124 ( .A(n119), .B(n105), .Y(n111) );
  NOR2X1 U125 ( .A(B[11]), .B(A[11]), .Y(n105) );
  NAND2X1 U126 ( .A(B[11]), .B(A[11]), .Y(n107) );
  OAI21X1 U127 ( .A(n112), .B(n123), .C(n109), .Y(n110) );
  XOR2X1 U128 ( .A(n113), .B(n123), .Y(SUM[10]) );
  OAI21X1 U129 ( .A(n124), .B(n30), .C(n31), .Y(n108) );
  NAND2X1 U130 ( .A(B[9]), .B(A[9]), .Y(n31) );
  NOR2X1 U131 ( .A(B[9]), .B(A[9]), .Y(n30) );
  OAI21X1 U132 ( .A(n34), .B(n114), .C(n33), .Y(n28) );
  NAND2X1 U133 ( .A(B[8]), .B(A[8]), .Y(n33) );
  NOR2X1 U134 ( .A(B[8]), .B(A[8]), .Y(n34) );
  NAND2X1 U135 ( .A(n121), .B(n109), .Y(n113) );
  NAND2X1 U136 ( .A(B[10]), .B(A[10]), .Y(n109) );
  NOR2X1 U137 ( .A(B[10]), .B(A[10]), .Y(n112) );
  INVX2 U3 ( .A(n93), .Y(n115) );
  INVX2 U4 ( .A(n99), .Y(n116) );
  INVX2 U5 ( .A(n101), .Y(n117) );
  INVX2 U6 ( .A(n104), .Y(n118) );
  INVX2 U7 ( .A(n107), .Y(n119) );
  INVX2 U8 ( .A(n109), .Y(n120) );
  INVX2 U9 ( .A(n112), .Y(n121) );
  INVX2 U10 ( .A(n31), .Y(n122) );
  INVX2 U11 ( .A(n108), .Y(n123) );
  INVX2 U12 ( .A(n28), .Y(n124) );
  INVX2 U13 ( .A(n34), .Y(n125) );
  INVX2 U14 ( .A(A[7]), .Y(n126) );
  INVX2 U15 ( .A(n37), .Y(n127) );
  INVX2 U16 ( .A(n43), .Y(n128) );
  INVX2 U17 ( .A(n45), .Y(n129) );
  INVX2 U18 ( .A(n51), .Y(n130) );
  INVX2 U19 ( .A(n53), .Y(n131) );
  INVX2 U20 ( .A(n59), .Y(n132) );
  INVX2 U21 ( .A(n61), .Y(n133) );
  INVX2 U22 ( .A(n67), .Y(n134) );
  INVX2 U23 ( .A(n69), .Y(n135) );
  INVX2 U24 ( .A(n75), .Y(n136) );
  INVX2 U25 ( .A(n77), .Y(n137) );
  INVX2 U26 ( .A(n83), .Y(n138) );
  INVX2 U27 ( .A(n85), .Y(n139) );
  INVX2 U28 ( .A(n91), .Y(n140) );
endmodule


module CannyEdge_DW02_mult_24 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[7][0] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][1] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[36] , \A1[35] , \A1[34] , \A1[33] ,
         \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] ,
         \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[4] ,
         \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n130, n131, n132, n133, n134, n135, n136,
         n137, n145, n143, n142, n141, n140, n139, n138, n13, n129, n114,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][30] , \SUMB[7][2] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][30] , \SUMB[6][2] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][30] , \SUMB[3][29] , \SUMB[3][28] ,
         \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] ,
         \SUMB[3][23] , \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] ,
         \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] , \SUMB[3][16] ,
         \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] ,
         \SUMB[3][11] , \SUMB[3][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][30] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[1][7] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][30] ,
         \CARRYB[7][2] , \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] ,
         \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] ,
         \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][1] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][30] , \CARRYB[6][2] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][30] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][30] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n144, n146, n147,
         n148, n149, n150, n151, n152, n153, n154;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n20), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n19), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n18), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n17), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n16), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n15), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  OR2X2 U5 ( .A(n116), .B(n109), .Y(n115) );
  OR2X2 U6 ( .A(n118), .B(n109), .Y(n117) );
  OR2X2 U7 ( .A(n120), .B(n109), .Y(n119) );
  OR2X2 U8 ( .A(n122), .B(n109), .Y(n121) );
  OR2X2 U9 ( .A(n124), .B(n109), .Y(n123) );
  OR2X2 U10 ( .A(n126), .B(n109), .Y(n125) );
  OR2X2 U11 ( .A(n128), .B(n109), .Y(n127) );
  AND2X1 U64 ( .A(\CARRYB[7][0] ), .B(\SUMB[7][1] ), .Y(n21) );
  NOR2X1 U65 ( .A(n111), .B(n115), .Y(n20) );
  NOR2X1 U66 ( .A(n112), .B(n117), .Y(n19) );
  NOR2X1 U67 ( .A(n113), .B(n119), .Y(n18) );
  NOR2X1 U68 ( .A(n144), .B(n121), .Y(n17) );
  NOR2X1 U69 ( .A(n146), .B(n123), .Y(n16) );
  NOR2X1 U70 ( .A(n147), .B(n125), .Y(n15) );
  NOR2X1 U71 ( .A(n148), .B(n127), .Y(n14) );
  NOR2X1 U75 ( .A(n154), .B(n148), .Y(\ab[7][7] ) );
  NOR2X1 U76 ( .A(n154), .B(n147), .Y(\ab[7][6] ) );
  NOR2X1 U77 ( .A(n154), .B(n146), .Y(\ab[7][5] ) );
  NOR2X1 U78 ( .A(n154), .B(n144), .Y(\ab[7][4] ) );
  NOR2X1 U79 ( .A(n154), .B(n113), .Y(\ab[7][3] ) );
  NOR2X1 U80 ( .A(n154), .B(n112), .Y(\ab[7][2] ) );
  NOR2X1 U81 ( .A(n154), .B(n111), .Y(\ab[7][1] ) );
  NOR2X1 U82 ( .A(n154), .B(n110), .Y(\ab[7][0] ) );
  NOR2X1 U83 ( .A(n153), .B(n148), .Y(\ab[6][7] ) );
  NOR2X1 U84 ( .A(n153), .B(n147), .Y(\ab[6][6] ) );
  NOR2X1 U85 ( .A(n153), .B(n146), .Y(\ab[6][5] ) );
  NOR2X1 U86 ( .A(n153), .B(n144), .Y(\ab[6][4] ) );
  NOR2X1 U87 ( .A(n153), .B(n113), .Y(\ab[6][3] ) );
  NOR2X1 U88 ( .A(n153), .B(n112), .Y(\ab[6][2] ) );
  NOR2X1 U89 ( .A(n153), .B(n111), .Y(\ab[6][1] ) );
  NOR2X1 U90 ( .A(n153), .B(n110), .Y(\ab[6][0] ) );
  NOR2X1 U91 ( .A(n152), .B(n148), .Y(\ab[5][7] ) );
  NOR2X1 U92 ( .A(n152), .B(n147), .Y(\ab[5][6] ) );
  NOR2X1 U93 ( .A(n152), .B(n146), .Y(\ab[5][5] ) );
  NOR2X1 U94 ( .A(n152), .B(n144), .Y(\ab[5][4] ) );
  NOR2X1 U95 ( .A(n152), .B(n113), .Y(\ab[5][3] ) );
  NOR2X1 U96 ( .A(n152), .B(n112), .Y(\ab[5][2] ) );
  NOR2X1 U97 ( .A(n152), .B(n111), .Y(\ab[5][1] ) );
  NOR2X1 U98 ( .A(n152), .B(n110), .Y(\ab[5][0] ) );
  NOR2X1 U99 ( .A(n151), .B(n148), .Y(\ab[4][7] ) );
  NOR2X1 U100 ( .A(n151), .B(n147), .Y(\ab[4][6] ) );
  NOR2X1 U101 ( .A(n151), .B(n146), .Y(\ab[4][5] ) );
  NOR2X1 U102 ( .A(n151), .B(n144), .Y(\ab[4][4] ) );
  NOR2X1 U103 ( .A(n151), .B(n113), .Y(\ab[4][3] ) );
  NOR2X1 U104 ( .A(n151), .B(n112), .Y(\ab[4][2] ) );
  NOR2X1 U105 ( .A(n151), .B(n111), .Y(\ab[4][1] ) );
  NOR2X1 U106 ( .A(n151), .B(n110), .Y(\ab[4][0] ) );
  NOR2X1 U107 ( .A(n150), .B(n148), .Y(\ab[3][7] ) );
  NOR2X1 U108 ( .A(n150), .B(n147), .Y(\ab[3][6] ) );
  NOR2X1 U109 ( .A(n150), .B(n146), .Y(\ab[3][5] ) );
  NOR2X1 U110 ( .A(n150), .B(n144), .Y(\ab[3][4] ) );
  NOR2X1 U111 ( .A(n150), .B(n113), .Y(\ab[3][3] ) );
  NOR2X1 U112 ( .A(n150), .B(n112), .Y(\ab[3][2] ) );
  NOR2X1 U113 ( .A(n150), .B(n111), .Y(\ab[3][1] ) );
  NOR2X1 U114 ( .A(n150), .B(n110), .Y(\ab[3][0] ) );
  NOR2X1 U115 ( .A(n149), .B(n148), .Y(\ab[2][7] ) );
  NOR2X1 U116 ( .A(n149), .B(n147), .Y(\ab[2][6] ) );
  NOR2X1 U117 ( .A(n149), .B(n146), .Y(\ab[2][5] ) );
  NOR2X1 U118 ( .A(n149), .B(n144), .Y(\ab[2][4] ) );
  NOR2X1 U119 ( .A(n149), .B(n113), .Y(\ab[2][3] ) );
  NOR2X1 U120 ( .A(n149), .B(n112), .Y(\ab[2][2] ) );
  NOR2X1 U121 ( .A(n149), .B(n111), .Y(\ab[2][1] ) );
  NOR2X1 U122 ( .A(n149), .B(n110), .Y(\ab[2][0] ) );
  NAND2X1 U124 ( .A(B[7]), .B(A[1]), .Y(n130) );
  XOR2X1 U125 ( .A(n128), .B(n131), .Y(\SUMB[1][6] ) );
  NAND2X1 U126 ( .A(B[7]), .B(A[0]), .Y(n131) );
  NAND2X1 U127 ( .A(B[6]), .B(A[1]), .Y(n128) );
  XOR2X1 U128 ( .A(n126), .B(n132), .Y(\SUMB[1][5] ) );
  NAND2X1 U129 ( .A(B[6]), .B(A[0]), .Y(n132) );
  NAND2X1 U130 ( .A(B[5]), .B(A[1]), .Y(n126) );
  XOR2X1 U131 ( .A(n124), .B(n133), .Y(\SUMB[1][4] ) );
  NAND2X1 U132 ( .A(B[5]), .B(A[0]), .Y(n133) );
  NAND2X1 U133 ( .A(B[4]), .B(A[1]), .Y(n124) );
  XOR2X1 U134 ( .A(n122), .B(n134), .Y(\SUMB[1][3] ) );
  NAND2X1 U135 ( .A(B[4]), .B(A[0]), .Y(n134) );
  NAND2X1 U136 ( .A(B[3]), .B(A[1]), .Y(n122) );
  XOR2X1 U137 ( .A(n120), .B(n135), .Y(\SUMB[1][2] ) );
  NAND2X1 U138 ( .A(B[3]), .B(A[0]), .Y(n135) );
  NAND2X1 U139 ( .A(B[2]), .B(A[1]), .Y(n120) );
  XOR2X1 U140 ( .A(n118), .B(n136), .Y(\SUMB[1][1] ) );
  NAND2X1 U141 ( .A(B[2]), .B(A[0]), .Y(n136) );
  NAND2X1 U142 ( .A(B[1]), .B(A[1]), .Y(n118) );
  XOR2X1 U146 ( .A(n116), .B(n137), .Y(PRODUCT[1]) );
  NAND2X1 U147 ( .A(B[1]), .B(A[0]), .Y(n137) );
  NAND2X1 U148 ( .A(B[0]), .B(A[1]), .Y(n116) );
  NOR2X1 U149 ( .A(n109), .B(n110), .Y(PRODUCT[0]) );
  XOR2X1 U153 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  CannyEdge_DW01_add_48 FS_1 ( .A({1'b0, \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \SUMB[7][0] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n3, 
        n4, n5, n6, n7, n8, n9, n10, n22, n30, n23, n31, n24, n32, n25, n33, 
        n26, n34, n27, n35, n28, n36, n29, n38, n37, n39, n40, n43, n41, n42, 
        n21, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  XOR2X1 U154 ( .A(\CARRYB[7][30] ), .B(n106), .Y(\A1[36] ) );
  AND2X1 U55 ( .A(n106), .B(\CARRYB[7][30] ), .Y(n3) );
  XOR2X1 U152 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  AND2X1 U41 ( .A(\CARRYB[7][1] ), .B(\SUMB[7][2] ), .Y(n42) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  XOR2X1 U151 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  AND2X1 U42 ( .A(\CARRYB[7][2] ), .B(\SUMB[7][3] ), .Y(n41) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  XOR2X1 U150 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  AND2X1 U40 ( .A(\CARRYB[7][3] ), .B(\SUMB[7][4] ), .Y(n43) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  XOR2X1 U181 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  AND2X1 U43 ( .A(\CARRYB[7][4] ), .B(\SUMB[7][5] ), .Y(n40) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  XOR2X1 U180 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  AND2X1 U45 ( .A(\CARRYB[7][5] ), .B(\SUMB[7][6] ), .Y(n39) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  XOR2X1 U179 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  AND2X1 U47 ( .A(\CARRYB[7][6] ), .B(\SUMB[7][7] ), .Y(n37) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n14), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U123 ( .A(n114), .B(n130), .Y(\SUMB[1][7] ) );
  XOR2X1 U175 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  AND2X1 U57 ( .A(\CARRYB[7][10] ), .B(\SUMB[7][11] ), .Y(n28) );
  XOR2X1 U174 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  AND2X1 U49 ( .A(\CARRYB[7][11] ), .B(\SUMB[7][12] ), .Y(n35) );
  FAX1 S4_11 ( .A(n106), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  XOR2X1 U171 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  AND2X1 U59 ( .A(\CARRYB[7][14] ), .B(\SUMB[7][15] ), .Y(n26) );
  XOR2X1 U170 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  AND2X1 U51 ( .A(\CARRYB[7][15] ), .B(\SUMB[7][16] ), .Y(n33) );
  FAX1 S4_15 ( .A(n106), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  XOR2X1 U167 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  AND2X1 U61 ( .A(\CARRYB[7][18] ), .B(\SUMB[7][19] ), .Y(n24) );
  XOR2X1 U166 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  AND2X1 U53 ( .A(\CARRYB[7][19] ), .B(\SUMB[7][20] ), .Y(n31) );
  FAX1 S4_19 ( .A(n106), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  XOR2X1 U163 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  AND2X1 U63 ( .A(\CARRYB[7][22] ), .B(\SUMB[7][23] ), .Y(n22) );
  XOR2X1 U162 ( .A(\SUMB[7][24] ), .B(\CARRYB[7][23] ), .Y(\A1[29] ) );
  AND2X1 U74 ( .A(\CARRYB[7][23] ), .B(\SUMB[7][24] ), .Y(n10) );
  FAX1 S4_23 ( .A(n106), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  XOR2X1 U159 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  AND2X1 U37 ( .A(\CARRYB[7][26] ), .B(\SUMB[7][27] ), .Y(n7) );
  XOR2X1 U158 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  AND2X1 U38 ( .A(\CARRYB[7][27] ), .B(\SUMB[7][28] ), .Y(n6) );
  FAX1 S4_27 ( .A(n106), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  XOR2X1 U178 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  AND2X1 U46 ( .A(\CARRYB[7][7] ), .B(\SUMB[7][8] ), .Y(n38) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n13), .C(n101), .YC(\CARRYB[2][7] ), .YS(
        \SUMB[2][7] ) );
  NOR2X1 U72 ( .A(n148), .B(n129), .Y(n13) );
  NAND2X1 U73 ( .A(n114), .B(A[1]), .Y(n129) );
  XOR2X1 U177 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  AND2X1 U56 ( .A(\CARRYB[7][8] ), .B(\SUMB[7][9] ), .Y(n29) );
  FAX1 S4_8 ( .A(n106), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S2_6_8 ( .A(n97), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_5_8 ( .A(n98), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_4_8 ( .A(n99), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_3_8 ( .A(n102), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_2_8 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][8] ), .YS(
        \SUMB[2][8] ) );
  XOR2X1 U157 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  AND2X1 U39 ( .A(\CARRYB[7][28] ), .B(\SUMB[7][29] ), .Y(n5) );
  FAX1 S4_28 ( .A(n106), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S2_6_28 ( .A(n97), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  XOR2X1 U161 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  AND2X1 U35 ( .A(\CARRYB[7][24] ), .B(\SUMB[7][25] ), .Y(n9) );
  FAX1 S4_24 ( .A(n106), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S2_6_24 ( .A(n97), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  XOR2X1 U165 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  AND2X1 U62 ( .A(\CARRYB[7][20] ), .B(\SUMB[7][21] ), .Y(n23) );
  FAX1 S4_20 ( .A(n106), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S2_6_20 ( .A(n97), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  XOR2X1 U169 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  AND2X1 U60 ( .A(\CARRYB[7][16] ), .B(\SUMB[7][17] ), .Y(n25) );
  FAX1 S4_16 ( .A(n106), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S2_6_16 ( .A(n97), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  XOR2X1 U173 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  AND2X1 U58 ( .A(\CARRYB[7][12] ), .B(\SUMB[7][13] ), .Y(n27) );
  FAX1 S4_12 ( .A(n106), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S2_6_12 ( .A(n97), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  XOR2X1 U176 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  AND2X1 U48 ( .A(\CARRYB[7][9] ), .B(\SUMB[7][10] ), .Y(n36) );
  FAX1 S4_10 ( .A(n106), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S2_6_11 ( .A(n97), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_5_12 ( .A(n98), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S4_9 ( .A(n106), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S2_6_10 ( .A(n97), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_5_11 ( .A(n98), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_4_12 ( .A(n99), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_6_9 ( .A(n97), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_5_10 ( .A(n98), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_4_11 ( .A(n99), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_3_12 ( .A(n102), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_5_9 ( .A(n98), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_4_10 ( .A(n99), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_3_11 ( .A(n102), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_2_12 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][12] ), .YS(
        \SUMB[2][12] ) );
  FAX1 S2_4_9 ( .A(n99), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_3_10 ( .A(n102), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_2_11 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][11] ), .YS(
        \SUMB[2][11] ) );
  FAX1 S2_3_9 ( .A(n102), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_2_10 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][10] ), .YS(
        \SUMB[2][10] ) );
  FAX1 S2_2_9 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][9] ), .YS(
        \SUMB[2][9] ) );
  XOR2X1 U172 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  AND2X1 U50 ( .A(\CARRYB[7][13] ), .B(\SUMB[7][14] ), .Y(n34) );
  FAX1 S4_14 ( .A(n106), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S2_6_15 ( .A(n97), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_5_16 ( .A(n98), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S4_13 ( .A(n106), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S2_6_14 ( .A(n97), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_5_15 ( .A(n98), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_4_16 ( .A(n99), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_6_13 ( .A(n97), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_5_14 ( .A(n98), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_4_15 ( .A(n99), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_3_16 ( .A(n102), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_5_13 ( .A(n98), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_4_14 ( .A(n99), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_3_15 ( .A(n102), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_2_16 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][16] ), .YS(
        \SUMB[2][16] ) );
  FAX1 S2_4_13 ( .A(n99), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_3_14 ( .A(n102), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_2_15 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][15] ), .YS(
        \SUMB[2][15] ) );
  FAX1 S2_3_13 ( .A(n102), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_2_14 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][14] ), .YS(
        \SUMB[2][14] ) );
  FAX1 S2_2_13 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][13] ), .YS(
        \SUMB[2][13] ) );
  XOR2X1 U168 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  AND2X1 U52 ( .A(\CARRYB[7][17] ), .B(\SUMB[7][18] ), .Y(n32) );
  FAX1 S4_18 ( .A(n106), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S2_6_19 ( .A(n97), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_5_20 ( .A(n98), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S4_17 ( .A(n106), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S2_6_18 ( .A(n97), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_5_19 ( .A(n98), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_4_20 ( .A(n99), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_6_17 ( .A(n97), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_5_18 ( .A(n98), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_4_19 ( .A(n99), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_3_20 ( .A(n102), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_5_17 ( .A(n98), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_4_18 ( .A(n99), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_3_19 ( .A(n102), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_2_20 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][20] ), .YS(
        \SUMB[2][20] ) );
  FAX1 S2_4_17 ( .A(n99), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_3_18 ( .A(n102), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_2_19 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][19] ), .YS(
        \SUMB[2][19] ) );
  FAX1 S2_3_17 ( .A(n102), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_2_18 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][18] ), .YS(
        \SUMB[2][18] ) );
  FAX1 S2_2_17 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][17] ), .YS(
        \SUMB[2][17] ) );
  XOR2X1 U164 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  AND2X1 U54 ( .A(\CARRYB[7][21] ), .B(\SUMB[7][22] ), .Y(n30) );
  FAX1 S4_22 ( .A(n106), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S2_6_23 ( .A(n97), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_5_24 ( .A(n98), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S4_21 ( .A(n106), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S2_6_22 ( .A(n97), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_5_23 ( .A(n98), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_4_24 ( .A(n99), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_6_21 ( .A(n97), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_5_22 ( .A(n98), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_4_23 ( .A(n99), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_3_24 ( .A(n102), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_5_21 ( .A(n98), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_4_22 ( .A(n99), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_3_23 ( .A(n102), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_2_24 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][24] ), .YS(
        \SUMB[2][24] ) );
  FAX1 S2_4_21 ( .A(n99), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_3_22 ( .A(n102), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_2_23 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][23] ), .YS(
        \SUMB[2][23] ) );
  FAX1 S2_3_21 ( .A(n102), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_2_22 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][22] ), .YS(
        \SUMB[2][22] ) );
  FAX1 S2_2_21 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][21] ), .YS(
        \SUMB[2][21] ) );
  XOR2X1 U160 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  AND2X1 U36 ( .A(\CARRYB[7][25] ), .B(\SUMB[7][26] ), .Y(n8) );
  FAX1 S4_26 ( .A(n106), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S2_6_27 ( .A(n97), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_5_28 ( .A(n98), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S4_25 ( .A(n106), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S2_6_26 ( .A(n97), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_5_27 ( .A(n98), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_4_28 ( .A(n99), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_6_25 ( .A(n97), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_5_26 ( .A(n98), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_4_27 ( .A(n99), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_3_28 ( .A(n102), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_5_25 ( .A(n98), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_4_26 ( .A(n99), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_3_27 ( .A(n102), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_2_28 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][28] ), .YS(
        \SUMB[2][28] ) );
  FAX1 S2_4_25 ( .A(n99), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_3_26 ( .A(n102), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_2_27 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][27] ), .YS(
        \SUMB[2][27] ) );
  FAX1 S2_3_25 ( .A(n102), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_2_26 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][26] ), .YS(
        \SUMB[2][26] ) );
  FAX1 S2_2_25 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][25] ), .YS(
        \SUMB[2][25] ) );
  XOR2X1 U156 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  AND2X1 U44 ( .A(\CARRYB[7][29] ), .B(\SUMB[7][30] ), .Y(n4) );
  FAX1 S5_30 ( .A(n106), .B(\CARRYB[6][30] ), .C(n97), .YC(\CARRYB[7][30] ), 
        .YS(\SUMB[7][30] ) );
  FAX1 S4_29 ( .A(n106), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S3_6_30 ( .A(n97), .B(\CARRYB[5][30] ), .C(n98), .YC(\CARRYB[6][30] ), 
        .YS(\SUMB[6][30] ) );
  FAX1 S2_6_29 ( .A(n97), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_5_30 ( .A(n98), .B(\CARRYB[4][30] ), .C(n99), .YC(\CARRYB[5][30] ), 
        .YS(\SUMB[5][30] ) );
  FAX1 S2_5_29 ( .A(n98), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_4_30 ( .A(n99), .B(\CARRYB[3][30] ), .C(n102), .YC(\CARRYB[4][30] ), 
        .YS(\SUMB[4][30] ) );
  FAX1 S2_4_29 ( .A(n99), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_3_30 ( .A(n102), .B(\CARRYB[2][30] ), .C(n103), .YC(\CARRYB[3][30] ), 
        .YS(\SUMB[3][30] ) );
  FAX1 S2_3_29 ( .A(n102), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_2_30 ( .A(n103), .B(n105), .C(n145), .YC(\CARRYB[2][30] ), .YS(
        \SUMB[2][30] ) );
  FAX1 S2_2_29 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][29] ), .YS(
        \SUMB[2][29] ) );
  NOR2X1 U145 ( .A(n109), .B(n107), .Y(n114) );
  AND2X1 U144 ( .A(A[1]), .B(B[9]), .Y(n145) );
  NOR2X1 U33 ( .A(n107), .B(n149), .Y(n143) );
  NOR2X1 U32 ( .A(n107), .B(n150), .Y(n142) );
  NOR2X1 U31 ( .A(n107), .B(n151), .Y(n141) );
  NOR2X1 U30 ( .A(n107), .B(n152), .Y(n140) );
  NOR2X1 U29 ( .A(n107), .B(n153), .Y(n139) );
  NOR2X1 U155 ( .A(n107), .B(n154), .Y(n138) );
  BUFX4 U12 ( .A(n139), .Y(n97) );
  BUFX4 U13 ( .A(n140), .Y(n98) );
  BUFX4 U14 ( .A(n141), .Y(n99) );
  XOR2X1 U15 ( .A(n108), .B(n145), .Y(n100) );
  INVX2 U16 ( .A(n100), .Y(n101) );
  BUFX4 U17 ( .A(n142), .Y(n102) );
  BUFX4 U18 ( .A(n143), .Y(n103) );
  NAND2X1 U19 ( .A(n145), .B(n114), .Y(n104) );
  INVX4 U20 ( .A(n104), .Y(n105) );
  BUFX4 U21 ( .A(n138), .Y(n106) );
  INVX2 U22 ( .A(B[9]), .Y(n107) );
  INVX2 U23 ( .A(n114), .Y(n108) );
  INVX2 U24 ( .A(A[0]), .Y(n109) );
  INVX2 U25 ( .A(B[0]), .Y(n110) );
  INVX2 U26 ( .A(B[1]), .Y(n111) );
  INVX2 U27 ( .A(B[2]), .Y(n112) );
  INVX2 U28 ( .A(B[3]), .Y(n113) );
  INVX2 U34 ( .A(B[4]), .Y(n144) );
  INVX2 U143 ( .A(B[5]), .Y(n146) );
  INVX2 U182 ( .A(B[6]), .Y(n147) );
  INVX2 U183 ( .A(B[7]), .Y(n148) );
  INVX2 U184 ( .A(A[2]), .Y(n149) );
  INVX2 U185 ( .A(A[3]), .Y(n150) );
  INVX2 U186 ( .A(A[4]), .Y(n151) );
  INVX2 U187 ( .A(A[5]), .Y(n152) );
  INVX2 U188 ( .A(A[6]), .Y(n153) );
  INVX2 U189 ( .A(A[7]), .Y(n154) );
endmodule


module CannyEdge ( dAddrRegRow, dAddrRegCol, bWE, bCE, InData, OutData, OPMode, 
        bOPEnable, dReadReg, dWriteReg, clk, rst_b );
  input [2:0] dAddrRegRow;
  input [2:0] dAddrRegCol;
  input [7:0] InData;
  output [7:0] OutData;
  input [2:0] OPMode;
  input [3:0] dReadReg;
  input [3:0] dWriteReg;
  input bWE, bCE, bOPEnable, clk, rst_b;
  wire   \regX[0][7] , \regX[0][6] , \regX[0][5] , \regX[0][4] , \regX[0][3] ,
         \regX[0][2] , \regX[0][1] , \regX[0][0] , \regX[1][7] , \regX[1][6] ,
         \regX[1][5] , \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] ,
         \regX[1][0] , \regX[3][7] , \regX[3][6] , \regX[3][5] , \regX[3][4] ,
         \regX[3][3] , \regX[3][2] , \regX[3][1] , \regX[3][0] , \regX[5][7] ,
         \regX[5][6] , \regX[5][5] , \regX[5][4] , \regX[5][3] , \regX[5][2] ,
         \regX[5][1] , \regX[5][0] , \regX[6][7] , \regX[6][6] , \regX[6][5] ,
         \regX[6][4] , \regX[6][3] , \regX[6][2] , \regX[6][1] , \regX[6][0] ,
         \regX[7][7] , \regX[7][6] , \regX[7][5] , \regX[7][4] , \regX[7][3] ,
         \regX[7][2] , \regX[7][1] , \regX[7][0] , \regX[8][7] , \regX[8][6] ,
         \regX[8][5] , \regX[8][4] , \regX[8][3] , \regX[8][2] , \regX[8][1] ,
         \regX[8][0] , \regX[9][7] , \regX[9][6] , \regX[9][5] , \regX[9][4] ,
         \regX[9][3] , \regX[9][2] , \regX[9][1] , \regX[9][0] , \regX[11][7] ,
         \regX[11][6] , \regX[11][5] , \regX[11][4] , \regX[11][3] ,
         \regX[11][2] , \regX[11][1] , \regX[11][0] , \regX[13][7] ,
         \regX[13][6] , \regX[13][5] , \regX[13][4] , \regX[13][3] ,
         \regX[13][2] , \regX[13][1] , \regX[13][0] , \regX[15][7] ,
         \regX[15][6] , \regX[15][5] , \regX[15][4] , \regX[15][3] ,
         \regX[15][2] , \regX[15][1] , \regX[15][0] , \regX[16][7] ,
         \regX[16][6] , \regX[16][5] , \regX[16][4] , \regX[16][3] ,
         \regX[16][2] , \regX[16][1] , \regX[16][0] , \regX[17][7] ,
         \regX[17][6] , \regX[17][5] , \regX[17][4] , \regX[17][3] ,
         \regX[17][2] , \regX[17][1] , \regX[17][0] , \regX[18][7] ,
         \regX[18][6] , \regX[18][5] , \regX[18][4] , \regX[18][3] ,
         \regX[18][2] , \regX[18][1] , \regX[18][0] , \regX[19][7] ,
         \regX[19][6] , \regX[19][5] , \regX[19][4] , \regX[19][3] ,
         \regX[19][2] , \regX[19][1] , \regX[19][0] , \regX[20][7] ,
         \regX[20][6] , \regX[20][5] , \regX[20][4] , \regX[20][3] ,
         \regX[20][2] , \regX[20][1] , \regX[20][0] , \regX[21][7] ,
         \regX[21][6] , \regX[21][5] , \regX[21][4] , \regX[21][3] ,
         \regX[21][2] , \regX[21][1] , \regX[21][0] , \regX[22][7] ,
         \regX[22][6] , \regX[22][5] , \regX[22][4] , \regX[22][3] ,
         \regX[22][2] , \regX[22][1] , \regX[22][0] , \regX[23][7] ,
         \regX[23][6] , \regX[23][5] , \regX[23][4] , \regX[23][3] ,
         \regX[23][2] , \regX[23][1] , \regX[23][0] , \regX[24][7] ,
         \regX[24][6] , \regX[24][5] , \regX[24][4] , \regX[24][3] ,
         \regX[24][2] , \regX[24][1] , \regX[24][0] , \regY[6][7] ,
         \regY[6][6] , \regY[6][5] , \regY[6][4] , \regY[6][3] , \regY[6][2] ,
         \regY[6][1] , \regY[6][0] , N971, N972, N973, N974, N975, N976, N977,
         N978, N979, N980, N981, N982, N983, \Out_bThres[0] , N1343, N1344,
         N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354,
         N1355, N1356, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382,
         N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1402, N1408, N1409, N1410, N1411, N1412,
         N1413, N1414, N1415, N1416, N1417, N1433, N1434, N1435, N1436, N1437,
         N1438, N1439, N1440, N1510, N1511, N1512, N1513, N1514, N1515, N1516,
         N1517, N1518, N1519, N1520, N1521, N1522, N1542, N1543, N1544, N1545,
         N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1570, N1571, N1572,
         N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582,
         N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1645, N1646,
         N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656,
         N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1707, N1708,
         N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1735, N1736,
         N1737, N1738, N1739, N1740, N1741, N1742, N1765, N1766, N1767, N1768,
         N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N2048, N2049,
         N2050, N2051, N2052, N2053, N2054, N2055, N2091, N2092, N2093, N2094,
         N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104,
         N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114,
         N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2155, N2156,
         N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166,
         N2167, N2168, N2169, N2170, N2171, N2236, N2237, N2238, N2239, N2240,
         N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250,
         N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260,
         N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270,
         N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280,
         N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290,
         N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300,
         N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310,
         N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320,
         N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330,
         N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340,
         N2341, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393,
         N2394, N2395, N2396, N2397, N2398, N2399, N2513, N2514, N2515, N2516,
         N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526,
         N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536,
         N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2549, N2558,
         N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568,
         N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2648, N2746,
         N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756,
         N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766,
         N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776,
         N2777, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832,
         N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2874,
         N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889,
         N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899,
         N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909,
         N2910, N2911, N2945, N3089, N3090, N3091, N3092, N3093, N3189, N3190,
         N3191, N3192, N3193, N3194, N3336, N3340, N3341, N3342, N3343, N3359,
         N3441, N3442, N3443, N3772, N3773, N3775, N3776, N3778, N3779, N3781,
         N3782, N3784, N3785, N3787, N3788, N3790, N3791, N3793, N3794, N3796,
         N3797, N3799, N3800, N3802, N3803, N3805, N3806, N3808, N3809, N3811,
         N3812, N3814, N3815, N3817, N3818, N3820, N3821, N3823, N3824, N3826,
         N3827, N3829, N3830, N3832, N3833, N3835, N3836, N3838, N3839, N3841,
         N3842, N3844, N3845, N3847, N3848, N3850, N3851, N3853, N3854, N3856,
         N3857, N3859, N3860, N3862, N3863, N3865, N3866, N3868, N3869, N3871,
         N3872, N3874, N3875, N3877, N3878, N3880, N3881, N3883, N3884, N3886,
         N3887, N3889, N3890, N3892, N3893, N3895, N3896, N3898, N3899, N3901,
         N3902, N3904, N3905, N3907, N3908, N3910, N3911, N3913, N3914, N3916,
         N3917, N3919, N3920, N3922, N3923, N3925, N3926, N3928, N3929, N3931,
         N3932, N3934, N3935, N3937, N3938, N3940, N3941, N3943, N3944, N3946,
         N3947, N3949, N3950, N3952, N3953, N3955, N3956, N3958, N3959, N3961,
         N3962, N3964, N3965, N3967, N3968, N3970, N3971, N3973, N3974, N3976,
         N3977, N3979, N3980, N3982, N3983, N3985, N3986, N3988, N3989, N3991,
         N3992, N3994, N3995, N3997, N3998, N4000, N4001, N4003, N4004, N4006,
         N4007, N4009, N4010, N4012, N4013, N4015, N4016, N4018, N4019, N4021,
         N4022, N4024, N4025, N4027, N4028, N4030, N4031, N4033, N4034, N4036,
         N4037, N4039, N4040, N4042, N4043, N4045, N4046, N4048, N4049, N4051,
         N4052, N4054, N4055, N4057, N4058, N4060, N4061, N4063, N4064, N4066,
         N4067, N4069, N4070, N4072, N4073, N4075, N4076, N4078, N4079, N4081,
         N4082, N4084, N4085, N4087, N4088, N4090, N4091, N4093, N4094, N4096,
         N4097, N4099, N4100, N4102, N4103, N4105, N4106, N4108, N4109, N4111,
         N4112, N4114, N4115, N4117, N4118, N4120, N4121, N4123, N4124, N4126,
         N4127, N4129, N4130, N4132, N4133, N4135, N4136, N4138, N4139, N4141,
         N4142, N4144, N4145, N4147, N4148, N4150, N4151, N4153, N4154, N4156,
         N4157, N4159, N4160, N4162, N4163, N4165, N4166, N4168, N4169, N4171,
         N4172, N4174, N4175, N4177, N4178, N4180, N4181, N4183, N4184, N4186,
         N4187, N4189, N4190, N4192, N4193, N4195, N4196, N4198, N4199, N4201,
         N4202, N4204, N4205, N4207, N4208, N4210, N4211, N4213, N4214, N4216,
         N4217, N4219, N4220, N4222, N4223, N4225, N4226, N4228, N4229, N4231,
         N4232, N4234, N4235, N4237, N4238, N4240, N4241, N4243, N4244, N4246,
         N4247, N4249, N4250, N4252, N4253, N4255, N4256, N4258, N4259, N4261,
         N4262, N4264, N4265, N4267, N4268, N4270, N4271, N4273, N4274, N4276,
         N4277, N4279, N4280, N4282, N4283, N4285, N4286, N4288, N4289, N4291,
         N4292, N4294, N4295, N4297, N4298, N4300, N4301, N4303, N4304, N4306,
         N4307, N4309, N4310, N4312, N4313, N4315, N4316, N4318, N4319, N4321,
         N4322, N4324, N4325, N4327, N4328, N4330, N4331, N4333, N4334, N4336,
         N4337, N4339, N4340, N4342, N4343, N4345, N4346, N4348, N4349, N4351,
         N4352, N4354, N4355, N4357, N4358, N4360, N4361, N4363, N4364, N4366,
         N4367, N4369, N4370, N4372, N4373, N4375, N4376, N4378, N4379, N4381,
         N4382, N4384, N4385, N4387, N4388, N4390, N4391, N4393, N4394, N4396,
         N4397, N4399, N4400, N4402, N4403, N4405, N4406, N4408, N4409, N4411,
         N4412, N4414, N4415, N4417, N4418, N4420, N4421, N4423, N4424, N4426,
         N4427, N4429, N4430, N4432, N4433, N4435, N4436, N4438, N4439, N4441,
         N4442, N4444, N4445, N4447, N4448, N4450, N4451, N4453, N4454, N4456,
         N4457, N4459, N4460, N4462, N4463, N4465, N4466, N4468, N4469, N4471,
         N4472, N4474, N4475, N4477, N4478, N4480, N4481, N4483, N4484, N4486,
         N4487, N4489, N4490, N4495, N4496, N4501, N4502, \U3/U63/Z_0 ,
         \U3/U63/Z_1 , \U3/U63/Z_2 , \U3/U63/Z_3 , \U3/U63/Z_4 , \U3/U63/Z_5 ,
         \U3/U63/Z_6 , \U3/U63/Z_7 , \U3/U64/Z_0 , \U3/U64/Z_1 , \U3/U64/Z_2 ,
         \U3/U64/Z_3 , \U3/U64/Z_4 , \U3/U64/Z_5 , \U3/U64/Z_6 , \U3/U64/Z_7 ,
         \U3/U65/Z_0 , \U3/U65/Z_1 , \U3/U65/Z_2 , \U3/U65/Z_3 , \U3/U65/Z_4 ,
         \U3/U65/Z_5 , \U3/U65/Z_6 , \U3/U65/Z_7 , \U3/U67/Z_1 , \U3/U68/Z_15 ,
         \U3/U68/Z_16 , \U3/U68/Z_17 , \U3/U68/Z_18 , \U3/U68/Z_19 ,
         \U3/U68/Z_20 , \U3/U68/Z_21 , \U3/U68/Z_22 , \U3/U68/Z_23 ,
         \U3/U68/Z_24 , \U3/U68/Z_25 , \U3/U68/Z_26 , \U3/U68/Z_27 ,
         \U3/U68/Z_28 , \U3/U68/Z_29 , \U3/U68/Z_30 , \U3/U68/Z_31 ,
         \U3/U69/Z_0 , \U3/U69/Z_1 , \U3/U69/Z_2 , \U3/U69/Z_3 , \U3/U69/Z_4 ,
         \U3/U69/Z_5 , \U3/U69/Z_6 , \U3/U69/Z_7 , \U3/U69/Z_8 , \U3/U69/Z_9 ,
         \U3/U69/Z_10 , \U3/U69/Z_11 , \U3/U69/Z_12 , \U3/U69/Z_13 ,
         \U3/U70/Z_0 , \U3/U70/Z_1 , \U3/U70/Z_2 , \U3/U70/Z_3 , \U3/U70/Z_4 ,
         \U3/U70/Z_5 , \U3/U70/Z_6 , \U3/U70/Z_7 , \U3/U70/Z_8 , \U3/U71/Z_15 ,
         \U3/U71/Z_16 , \U3/U71/Z_17 , \U3/U71/Z_18 , \U3/U71/Z_19 ,
         \U3/U71/Z_20 , \U3/U71/Z_21 , \U3/U71/Z_22 , \U3/U71/Z_23 ,
         \U3/U71/Z_24 , \U3/U71/Z_25 , \U3/U71/Z_26 , \U3/U71/Z_27 ,
         \U3/U71/Z_28 , \U3/U71/Z_29 , \U3/U71/Z_30 , \U3/U71/Z_31 ,
         \U3/U72/Z_15 , \U3/U72/Z_16 , \U3/U72/Z_17 , \U3/U72/Z_18 ,
         \U3/U72/Z_19 , \U3/U72/Z_20 , \U3/U72/Z_21 , \U3/U72/Z_22 ,
         \U3/U72/Z_23 , \U3/U72/Z_24 , \U3/U72/Z_25 , \U3/U72/Z_26 ,
         \U3/U72/Z_27 , \U3/U72/Z_28 , \U3/U72/Z_29 , \U3/U72/Z_30 ,
         \U3/U72/Z_31 , \U3/U73/Z_15 , \U3/U73/Z_16 , \U3/U73/Z_17 ,
         \U3/U73/Z_18 , \U3/U73/Z_19 , \U3/U73/Z_20 , \U3/U73/Z_21 ,
         \U3/U73/Z_22 , \U3/U73/Z_23 , \U3/U73/Z_24 , \U3/U73/Z_25 ,
         \U3/U73/Z_26 , \U3/U73/Z_27 , \U3/U73/Z_28 , \U3/U73/Z_29 ,
         \U3/U73/Z_30 , \U3/U73/Z_31 , \U3/U74/Z_15 , \U3/U74/Z_16 ,
         \U3/U74/Z_17 , \U3/U74/Z_18 , \U3/U74/Z_19 , \U3/U74/Z_20 ,
         \U3/U74/Z_21 , \U3/U74/Z_22 , \U3/U74/Z_23 , \U3/U74/Z_24 ,
         \U3/U74/Z_25 , \U3/U74/Z_26 , \U3/U74/Z_27 , \U3/U74/Z_28 ,
         \U3/U74/Z_29 , \U3/U74/Z_30 , \U3/U74/Z_31 , \U3/U75/Z_0 ,
         \U3/U75/Z_1 , \U3/U75/Z_2 , \U3/U75/Z_3 , \U3/U75/Z_4 , \U3/U75/Z_5 ,
         \U3/U75/Z_6 , \U3/U75/Z_7 , \U3/U75/Z_8 , \U3/U75/Z_9 , \U3/U75/Z_10 ,
         \U3/U75/Z_11 , \U3/U75/Z_12 , \U3/U75/Z_13 , \U3/U75/Z_14 ,
         \U3/U76/Z_10 , \U3/U76/Z_11 , \U3/U76/Z_12 , \U3/U76/Z_13 ,
         \U3/U76/Z_14 , \U3/U77/Z_15 , \U3/U77/Z_16 , \U3/U77/Z_17 ,
         \U3/U77/Z_18 , \U3/U77/Z_19 , \U3/U77/Z_20 , \U3/U77/Z_21 ,
         \U3/U77/Z_22 , \U3/U77/Z_23 , \U3/U77/Z_24 , \U3/U77/Z_25 ,
         \U3/U77/Z_26 , \U3/U77/Z_27 , \U3/U77/Z_28 , \U3/U77/Z_29 ,
         \U3/U77/Z_30 , \U3/U77/Z_31 , \U3/U77/DATA2_15 , \U3/U77/DATA2_16 ,
         \U3/U77/DATA2_17 , \U3/U77/DATA2_18 , \U3/U77/DATA2_19 ,
         \U3/U77/DATA2_20 , \U3/U77/DATA2_21 , \U3/U77/DATA2_22 ,
         \U3/U77/DATA2_23 , \U3/U77/DATA2_24 , \U3/U77/DATA2_25 ,
         \U3/U77/DATA2_26 , \U3/U77/DATA2_27 , \U3/U77/DATA2_28 ,
         \U3/U77/DATA2_29 , \U3/U77/DATA2_30 , \U3/U77/DATA2_31 , \U3/U78/Z_0 ,
         \U3/U78/Z_1 , \U3/U78/Z_2 , \U3/U78/Z_3 , \U3/U78/Z_4 , \U3/U78/Z_5 ,
         \U3/U78/Z_6 , \U3/U78/Z_7 , \U3/U78/Z_8 , \U3/U78/Z_9 , \U3/U78/Z_10 ,
         \U3/U78/Z_11 , \U3/U78/Z_12 , \U3/U78/Z_13 , \U3/U78/Z_14 ,
         \U3/U78/Z_15 , \U3/U78/Z_16 , \U3/U78/Z_17 , \U3/U78/Z_18 ,
         \U3/U78/Z_19 , \U3/U78/Z_20 , \U3/U78/Z_21 , \U3/U78/Z_22 ,
         \U3/U78/Z_23 , \U3/U78/Z_24 , \U3/U78/Z_25 , \U3/U78/Z_26 ,
         \U3/U78/Z_27 , \U3/U78/Z_28 , \U3/U78/Z_29 , \U3/U78/Z_30 ,
         \U3/U78/Z_31 , \U3/U79/Z_0 , \U3/U79/Z_1 , \U3/U79/Z_2 , \U3/U79/Z_3 ,
         \U3/U79/Z_4 , \U3/U79/Z_5 , \U3/U79/Z_6 , \U3/U79/Z_7 , \U3/U79/Z_8 ,
         \U3/U79/Z_9 , \U3/U79/Z_10 , \U3/U79/Z_11 , \U3/U79/Z_12 ,
         \U3/U79/Z_13 , \U3/U79/Z_14 , \U3/U79/Z_15 , \U3/U79/Z_16 ,
         \U3/U79/Z_17 , \U3/U79/Z_18 , \U3/U79/Z_19 , \U3/U79/Z_20 ,
         \U3/U79/Z_21 , \U3/U79/Z_22 , \U3/U79/Z_23 , \U3/U79/Z_24 ,
         \U3/U79/Z_25 , \U3/U79/Z_26 , \U3/U79/Z_27 , \U3/U79/Z_28 ,
         \U3/U79/Z_29 , \U3/U79/Z_30 , \U3/U79/Z_31 , \U3/U81/Z_0 ,
         \U3/U81/Z_1 , \U3/U81/Z_2 , \U3/U81/Z_3 , \U3/U81/Z_4 , \U3/U81/Z_5 ,
         \U3/U81/Z_6 , \U3/U81/Z_7 , \U3/U82/Z_0 , \U3/U82/Z_1 , \U3/U82/Z_2 ,
         \U3/U82/Z_3 , \U3/U82/Z_4 , \U3/U82/Z_5 , \U3/U82/Z_6 , \U3/U82/Z_7 ,
         \U3/U82/Z_8 , \U3/U82/Z_9 , \U3/U82/Z_10 , \U3/U82/Z_11 ,
         \U3/U82/Z_12 , \U3/U82/Z_13 , \U3/U82/Z_14 , \U3/U82/Z_15 ,
         \U3/U82/Z_16 , \U3/U82/Z_17 , \U3/U82/Z_18 , \U3/U82/Z_19 ,
         \U3/U82/Z_20 , \U3/U82/Z_21 , \U3/U82/Z_22 , \U3/U82/Z_23 ,
         \U3/U82/Z_24 , \U3/U82/Z_25 , \U3/U82/Z_26 , \U3/U82/Z_27 ,
         \U3/U82/Z_28 , \U3/U82/Z_29 , \U3/U82/Z_30 , \U3/U82/Z_31 ,
         \U3/U84/Z_0 , \U3/U84/Z_1 , \U3/U84/Z_2 , \U3/U84/Z_3 , \U3/U84/Z_4 ,
         \U3/U84/Z_5 , \U3/U84/Z_6 , \U3/U84/Z_7 , \U3/U85/Z_0 , \U3/U85/Z_1 ,
         \U3/U85/Z_2 , \U3/U85/Z_3 , \U3/U85/Z_4 , \U3/U85/Z_5 , \U3/U85/Z_6 ,
         \U3/U85/Z_7 , \U3/U85/Z_8 , \U3/U85/Z_9 , \U3/U85/Z_10 ,
         \U3/U85/Z_11 , \U3/U85/Z_12 , \U3/U85/Z_13 , \U3/U85/Z_14 ,
         \U3/U85/Z_15 , \U3/U85/Z_16 , \U3/U85/Z_17 , \U3/U85/Z_18 ,
         \U3/U85/Z_19 , \U3/U85/Z_20 , \U3/U85/Z_21 , \U3/U85/Z_22 ,
         \U3/U85/Z_23 , \U3/U85/Z_24 , \U3/U85/Z_25 , \U3/U85/Z_26 ,
         \U3/U85/Z_27 , \U3/U85/Z_28 , \U3/U85/Z_29 , \U3/U85/Z_30 ,
         \U3/U85/Z_31 , \U3/U87/Z_0 , \U3/U87/Z_1 , \U3/U87/Z_2 , \U3/U87/Z_3 ,
         \U3/U87/Z_4 , \U3/U87/Z_5 , \U3/U87/Z_6 , \U3/U87/Z_7 , \U3/U88/Z_0 ,
         \U3/U88/Z_1 , \U3/U88/Z_2 , \U3/U88/Z_3 , \U3/U88/Z_4 , \U3/U88/Z_5 ,
         \U3/U88/Z_6 , \U3/U88/Z_7 , \U3/U88/Z_8 , \U3/U88/Z_9 , \U3/U88/Z_10 ,
         \U3/U88/Z_11 , \U3/U88/Z_12 , \U3/U88/Z_13 , \U3/U88/Z_14 ,
         \U3/U88/Z_15 , \U3/U88/Z_16 , \U3/U88/Z_17 , \U3/U88/Z_18 ,
         \U3/U88/Z_19 , \U3/U88/Z_20 , \U3/U88/Z_21 , \U3/U88/Z_22 ,
         \U3/U88/Z_23 , \U3/U88/Z_24 , \U3/U88/Z_25 , \U3/U88/Z_26 ,
         \U3/U88/Z_27 , \U3/U88/Z_28 , \U3/U88/Z_29 , \U3/U88/Z_30 ,
         \U3/U90/Z_0 , \U3/U91/Z_0 , \U3/U91/Z_1 , \U3/U91/Z_2 , \U3/U91/Z_3 ,
         \U3/U91/Z_4 , \U3/U91/Z_5 , \U3/U91/Z_6 , \U3/U91/Z_7 , \U3/U93/Z_0 ,
         \U3/U93/Z_1 , \U3/U93/Z_2 , \U3/U93/Z_3 , \U3/U93/Z_4 , \U3/U93/Z_5 ,
         \U3/U93/Z_6 , \U3/U93/Z_7 , \U3/U93/Z_8 , \U3/U93/Z_9 , \U3/U93/Z_10 ,
         \U3/U93/Z_11 , \U3/U93/Z_12 , \U3/U93/Z_13 , \U3/U93/Z_14 ,
         \U3/U93/Z_15 , \U3/U93/Z_16 , \U3/U93/Z_17 , \U3/U93/Z_18 ,
         \U3/U93/Z_19 , \U3/U93/Z_20 , \U3/U93/Z_21 , \U3/U93/Z_22 ,
         \U3/U93/Z_23 , \U3/U93/Z_24 , \U3/U93/Z_25 , \U3/U93/Z_26 ,
         \U3/U93/Z_27 , \U3/U93/Z_28 , \U3/U93/Z_29 , \U3/U93/Z_30 ,
         \U3/U93/Z_31 , \U3/U94/Z_0 , \U3/U94/Z_1 , \U3/U94/Z_2 , \U3/U94/Z_3 ,
         \U3/U94/Z_4 , \U3/U94/Z_5 , \U3/U94/Z_6 , \U3/U94/Z_7 , \U3/U94/Z_8 ,
         \U3/U94/Z_9 , \U3/U94/Z_10 , \U3/U94/Z_11 , \U3/U94/Z_12 ,
         \U3/U94/Z_13 , \U3/U94/Z_14 , \U3/U94/Z_15 , \U3/U94/Z_16 ,
         \U3/U94/Z_17 , \U3/U94/Z_18 , \U3/U94/Z_19 , \U3/U94/Z_20 ,
         \U3/U94/Z_21 , \U3/U94/Z_22 , \U3/U94/Z_23 , \U3/U94/Z_24 ,
         \U3/U94/Z_25 , \U3/U94/Z_26 , \U3/U94/Z_27 , \U3/U94/Z_28 ,
         \U3/U94/Z_29 , \U3/U94/Z_31 , \U3/U95/Z_0 , \U3/U96/Z_0 ,
         \U3/U97/Z_0 , \U3/U98/Z_0 , \U3/U98/Z_1 , \U3/U98/Z_2 , \U3/U98/Z_3 ,
         \U3/U98/Z_4 , \U3/U98/Z_5 , \U3/U98/Z_6 , \U3/U98/Z_7 , \U3/U100/Z_0 ,
         \U3/U100/Z_1 , \U3/U100/Z_2 , \U3/U100/Z_3 , \U3/U100/Z_4 ,
         \U3/U100/Z_6 , \U3/U101/Z_0 , \U3/U101/Z_1 , \U3/U101/Z_2 ,
         \U3/U101/Z_3 , \U3/U101/Z_6 , \U3/U105/Z_0 , \U3/U105/Z_1 ,
         \U3/U105/Z_2 , \U3/U105/Z_3 , \U3/U106/Z_1 , \U3/U106/Z_3 ,
         \U3/U107/Z_0 , \U3/U109/Z_2 , \U3/U110/Z_1 , \U3/U110/Z_2 ,
         \U3/U110/Z_3 , \U3/U110/Z_4 , \U3/U110/Z_5 , \U3/U110/Z_6 ,
         \U3/U110/Z_7 , \U3/U118/Z_0 , \U3/U118/Z_1 , \U3/U118/Z_2 ,
         \U3/U118/Z_3 , \U3/U118/Z_4 , \U3/U118/Z_5 , \U3/U118/Z_6 ,
         \U3/U118/Z_7 , \U3/U118/Z_8 , \U3/U118/Z_9 , \U3/U118/Z_10 ,
         \U3/U118/Z_11 , \U3/U118/Z_12 , \U3/U118/Z_13 , \U3/U118/Z_14 ,
         \U3/U118/Z_15 , \U3/U118/Z_16 , \U3/U118/Z_17 , \U3/U118/Z_18 ,
         \U3/U118/Z_19 , \U3/U118/Z_20 , \U3/U118/Z_21 , \U3/U118/Z_22 ,
         \U3/U118/Z_23 , \U3/U118/Z_24 , \U3/U118/Z_25 , \U3/U118/Z_26 ,
         \U3/U118/Z_27 , \U3/U118/Z_28 , \U3/U118/Z_29 , \U3/U118/Z_30 ,
         \U3/U118/Z_31 , \U3/U119/Z_0 , \U3/U119/Z_1 , \U3/U119/Z_2 ,
         \U3/U119/Z_3 , \U3/U119/Z_4 , \U3/U119/Z_5 , \U3/U119/Z_6 ,
         \U3/U119/Z_7 , \U3/U119/Z_8 , \U3/U119/Z_9 , \U3/U119/Z_10 ,
         \U3/U119/Z_11 , \U3/U119/Z_12 , \U3/U119/Z_13 , \U3/U119/Z_14 ,
         \U3/U119/Z_15 , \U3/U119/Z_16 , \U3/U119/Z_17 , \U3/U119/Z_18 ,
         \U3/U119/Z_19 , \U3/U119/Z_20 , \U3/U119/Z_21 , \U3/U119/Z_22 ,
         \U3/U119/Z_23 , \U3/U119/Z_24 , \U3/U119/Z_25 , \U3/U119/Z_26 ,
         \U3/U119/Z_27 , \U3/U119/Z_28 , \U3/U119/Z_29 , \U3/U119/Z_31 ,
         \U3/U121/Z_0 , \U3/U121/Z_1 , \U3/U121/Z_2 , \U3/U121/Z_3 ,
         \U3/U121/Z_4 , \U3/U121/Z_5 , \U3/U121/Z_6 , \U3/U121/Z_7 ,
         \U3/U122/Z_0 , \U3/U122/Z_1 , \U3/U122/Z_2 , \U3/U122/Z_3 ,
         \U3/U122/Z_4 , \U3/U122/Z_5 , \U3/U122/Z_6 , \U3/U122/Z_7 ,
         \U3/U122/Z_8 , \U3/U122/Z_9 , \U3/U122/Z_10 , \U3/U122/Z_11 ,
         \U3/U122/Z_12 , \U3/U122/Z_13 , \U3/U122/Z_14 , \U3/U122/Z_15 ,
         \U3/U122/Z_16 , \U3/U122/Z_17 , \U3/U122/Z_18 , \U3/U122/Z_19 ,
         \U3/U122/Z_20 , \U3/U122/Z_21 , \U3/U122/Z_22 , \U3/U122/Z_23 ,
         \U3/U122/Z_24 , \U3/U122/Z_25 , \U3/U122/Z_26 , \U3/U122/Z_27 ,
         \U3/U122/Z_28 , \U3/U122/Z_29 , \U3/U124/Z_0 , \U3/U125/Z_0 ,
         \U3/U125/Z_1 , \U3/U125/Z_2 , \U3/U125/Z_3 , \U3/U125/Z_4 ,
         \U3/U125/Z_5 , \U3/U125/Z_6 , \U3/U125/Z_7 , \U3/U134/Z_0 ,
         \U3/U134/Z_1 , \U3/U134/Z_2 , \U3/U134/Z_3 , \U3/U134/Z_4 ,
         \U3/U134/Z_5 , \U3/U134/Z_6 , \U3/U134/Z_7 , \U3/U134/Z_8 ,
         \U3/U134/Z_9 , \U3/U134/Z_10 , \U3/U136/Z_0 , n4565, n4567, n4569,
         n4571, n4573, n4575, n4577, n4579, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5396, n5397, n5398, n5409, n8287, n8288, n8289,
         n8291, n8303, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815,
         N2814, N2813, N2812, N2811, N2810, N2481, N2480, N2479, N2478, N2477,
         N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467,
         N2466, N2465, N2464, N2417, N2416, N2415, N2414, N2413, N2412, N2411,
         N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401,
         N2400, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195,
         N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185,
         N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175,
         N2174, N2173, N2172, N2154, N2153, N2152, N2151, N2150, N2149, N2148,
         N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138,
         N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128,
         N2127, N2126, N2125, N2124, N2123, N2090, N2089, N2088, N2087, N2086,
         N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076,
         N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023,
         N2022, N2021, N2020, N2019, N2018, N2002, N2001, N2000, N1999, N1998,
         N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988,
         N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963,
         N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953,
         N1952, N1951, N1950, N1949, N1942, N1941, N1940, N1939, N1938, N1937,
         N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927,
         N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1912,
         N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902,
         N1901, N1900, N1899, N1898, N1896, N1895, N1894, N1893, N1892, N1891,
         N1890, N1889, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875,
         N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865,
         N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1852, N1851, N1850,
         N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840,
         N1839, N1838, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829,
         N1828, N1827, N1826, N1825, N1824, N1822, N1821, N1820, N1819, N1818,
         N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1806,
         N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796,
         N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786,
         N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1762, N1761,
         N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751,
         N1750, N1749, N1748, N1732, N1731, N1730, N1729, N1728, N1727, N1726,
         N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1672, N1671,
         N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661,
         N1660, N1659, N1658, N1642, N1641, N1640, N1639, N1638, N1637, N1636,
         N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1612, N1611,
         N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601,
         N1600, N1599, N1598, N1596, N1595, N1594, N1593, N1592, N1591, N1590,
         N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1569, N1568, N1566,
         N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556,
         N1555, N1554, N1553, N1541, N1540, N1539, N1536, N1535, N1534, N1533,
         N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1509,
         N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497,
         N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487,
         N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1462,
         N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452,
         N1451, N1450, N1449, N1448, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853;
  wire   [7:0] Out_gf;
  wire   [1:0] IntSignal;
  wire   [14:7] tpSum;
  wire   [31:0] Gx;
  wire   [31:0] Gy;
  tri   [7:0] OutData;
  tri   [31:0] fGy;
  tri   [31:0] fGx;
  tri   [1:0] dx;
  tri   [1:0] dy;
  tri   \regZ[0][7] ;
  tri   \regZ[0][6] ;
  tri   \regZ[0][5] ;
  tri   \regZ[0][4] ;
  tri   \regZ[0][3] ;
  tri   \regZ[0][2] ;
  tri   \regZ[0][1] ;
  tri   \regZ[0][0] ;
  tri   \regZ[1][7] ;
  tri   \regZ[1][6] ;
  tri   \regZ[1][5] ;
  tri   \regZ[1][4] ;
  tri   \regZ[1][3] ;
  tri   \regZ[1][2] ;
  tri   \regZ[1][1] ;
  tri   \regZ[1][0] ;
  tri   \regZ[2][7] ;
  tri   \regZ[2][6] ;
  tri   \regZ[2][5] ;
  tri   \regZ[2][4] ;
  tri   \regZ[2][3] ;
  tri   \regZ[2][2] ;
  tri   \regZ[2][1] ;
  tri   \regZ[2][0] ;
  tri   \regZ[3][7] ;
  tri   \regZ[3][6] ;
  tri   \regZ[3][5] ;
  tri   \regZ[3][4] ;
  tri   \regZ[3][3] ;
  tri   \regZ[3][2] ;
  tri   \regZ[3][1] ;
  tri   \regZ[3][0] ;
  tri   \regZ[4][7] ;
  tri   \regZ[4][6] ;
  tri   \regZ[4][5] ;
  tri   \regZ[4][4] ;
  tri   \regZ[4][3] ;
  tri   \regZ[4][2] ;
  tri   \regZ[4][1] ;
  tri   \regZ[4][0] ;
  tri   \regZ[5][7] ;
  tri   \regZ[5][6] ;
  tri   \regZ[5][5] ;
  tri   \regZ[5][4] ;
  tri   \regZ[5][3] ;
  tri   \regZ[5][2] ;
  tri   \regZ[5][1] ;
  tri   \regZ[5][0] ;
  tri   \regZ[6][7] ;
  tri   \regZ[6][6] ;
  tri   \regZ[6][5] ;
  tri   \regZ[6][4] ;
  tri   \regZ[6][3] ;
  tri   \regZ[6][2] ;
  tri   \regZ[6][1] ;
  tri   \regZ[6][0] ;
  tri   \regZ[7][7] ;
  tri   \regZ[7][6] ;
  tri   \regZ[7][5] ;
  tri   \regZ[7][4] ;
  tri   \regZ[7][3] ;
  tri   \regZ[7][2] ;
  tri   \regZ[7][1] ;
  tri   \regZ[7][0] ;
  tri   \regZ[8][7] ;
  tri   \regZ[8][6] ;
  tri   \regZ[8][5] ;
  tri   \regZ[8][4] ;
  tri   \regZ[8][3] ;
  tri   \regZ[8][2] ;
  tri   \regZ[8][1] ;
  tri   \regZ[8][0] ;
  tri   \regZ[9][7] ;
  tri   \regZ[9][6] ;
  tri   \regZ[9][5] ;
  tri   \regZ[9][4] ;
  tri   \regZ[9][3] ;
  tri   \regZ[9][2] ;
  tri   \regZ[9][1] ;
  tri   \regZ[9][0] ;
  tri   \regZ[10][7] ;
  tri   \regZ[10][6] ;
  tri   \regZ[10][5] ;
  tri   \regZ[10][4] ;
  tri   \regZ[10][3] ;
  tri   \regZ[10][2] ;
  tri   \regZ[10][1] ;
  tri   \regZ[10][0] ;
  tri   \regZ[11][7] ;
  tri   \regZ[11][6] ;
  tri   \regZ[11][5] ;
  tri   \regZ[11][4] ;
  tri   \regZ[11][3] ;
  tri   \regZ[11][2] ;
  tri   \regZ[11][1] ;
  tri   \regZ[11][0] ;
  tri   \regZ[12][7] ;
  tri   \regZ[12][6] ;
  tri   \regZ[12][5] ;
  tri   \regZ[12][4] ;
  tri   \regZ[12][3] ;
  tri   \regZ[12][2] ;
  tri   \regZ[12][1] ;
  tri   \regZ[12][0] ;
  tri   \regZ[13][7] ;
  tri   \regZ[13][6] ;
  tri   \regZ[13][5] ;
  tri   \regZ[13][4] ;
  tri   \regZ[13][3] ;
  tri   \regZ[13][2] ;
  tri   \regZ[13][1] ;
  tri   \regZ[13][0] ;
  tri   \regZ[14][7] ;
  tri   \regZ[14][6] ;
  tri   \regZ[14][5] ;
  tri   \regZ[14][4] ;
  tri   \regZ[14][3] ;
  tri   \regZ[14][2] ;
  tri   \regZ[14][1] ;
  tri   \regZ[14][0] ;
  tri   \regZ[15][7] ;
  tri   \regZ[15][6] ;
  tri   \regZ[15][5] ;
  tri   \regZ[15][4] ;
  tri   \regZ[15][3] ;
  tri   \regZ[15][2] ;
  tri   \regZ[15][1] ;
  tri   \regZ[15][0] ;
  tri   \regZ[16][7] ;
  tri   \regZ[16][6] ;
  tri   \regZ[16][5] ;
  tri   \regZ[16][4] ;
  tri   \regZ[16][3] ;
  tri   \regZ[16][2] ;
  tri   \regZ[16][1] ;
  tri   \regZ[16][0] ;
  tri   \regZ[17][7] ;
  tri   \regZ[17][6] ;
  tri   \regZ[17][5] ;
  tri   \regZ[17][4] ;
  tri   \regZ[17][3] ;
  tri   \regZ[17][2] ;
  tri   \regZ[17][1] ;
  tri   \regZ[17][0] ;
  tri   \regZ[18][7] ;
  tri   \regZ[18][6] ;
  tri   \regZ[18][5] ;
  tri   \regZ[18][4] ;
  tri   \regZ[18][3] ;
  tri   \regZ[18][2] ;
  tri   \regZ[18][1] ;
  tri   \regZ[18][0] ;
  tri   \regZ[19][7] ;
  tri   \regZ[19][6] ;
  tri   \regZ[19][5] ;
  tri   \regZ[19][4] ;
  tri   \regZ[19][3] ;
  tri   \regZ[19][2] ;
  tri   \regZ[19][1] ;
  tri   \regZ[19][0] ;
  tri   \regZ[20][7] ;
  tri   \regZ[20][6] ;
  tri   \regZ[20][5] ;
  tri   \regZ[20][4] ;
  tri   \regZ[20][3] ;
  tri   \regZ[20][2] ;
  tri   \regZ[20][1] ;
  tri   \regZ[20][0] ;
  tri   \regZ[21][7] ;
  tri   \regZ[21][6] ;
  tri   \regZ[21][5] ;
  tri   \regZ[21][4] ;
  tri   \regZ[21][3] ;
  tri   \regZ[21][2] ;
  tri   \regZ[21][1] ;
  tri   \regZ[21][0] ;
  tri   \regZ[22][7] ;
  tri   \regZ[22][6] ;
  tri   \regZ[22][5] ;
  tri   \regZ[22][4] ;
  tri   \regZ[22][3] ;
  tri   \regZ[22][2] ;
  tri   \regZ[22][1] ;
  tri   \regZ[22][0] ;
  tri   \regZ[23][7] ;
  tri   \regZ[23][6] ;
  tri   \regZ[23][5] ;
  tri   \regZ[23][4] ;
  tri   \regZ[23][3] ;
  tri   \regZ[23][2] ;
  tri   \regZ[23][1] ;
  tri   \regZ[23][0] ;
  tri   \regZ[24][7] ;
  tri   \regZ[24][6] ;
  tri   \regZ[24][5] ;
  tri   \regZ[24][4] ;
  tri   \regZ[24][3] ;
  tri   \regZ[24][2] ;
  tri   \regZ[24][1] ;
  tri   \regZ[24][0] ;
  tri   [7:0] Out_gradient;
  tri   [7:0] Out_direction;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80;

  DFFPOSX1 \OutData_tri_enable_reg[7]  ( .D(n5389), .CLK(clk), .Q(N4469) );
  DFFPOSX1 \OutData_tri_enable_reg[6]  ( .D(n5388), .CLK(clk), .Q(N4472) );
  DFFPOSX1 \OutData_tri_enable_reg[5]  ( .D(n5387), .CLK(clk), .Q(N4475) );
  DFFPOSX1 \OutData_tri_enable_reg[4]  ( .D(n5386), .CLK(clk), .Q(N4478) );
  DFFPOSX1 \OutData_tri_enable_reg[3]  ( .D(n5385), .CLK(clk), .Q(N4481) );
  DFFPOSX1 \OutData_tri_enable_reg[2]  ( .D(n5384), .CLK(clk), .Q(N4484) );
  DFFPOSX1 \OutData_tri_enable_reg[1]  ( .D(n5383), .CLK(clk), .Q(N4487) );
  DFFPOSX1 \OutData_tri_enable_reg[0]  ( .D(n5382), .CLK(clk), .Q(N4490) );
  DFFSR \IntSignal_reg[0]  ( .D(n5381), .CLK(clk), .R(rst_b), .S(rst_b), .Q(
        IntSignal[0]) );
  DFFSR \IntSignal_reg[1]  ( .D(n15368), .CLK(clk), .R(rst_b), .S(rst_b), .Q(
        IntSignal[1]) );
  DFFPOSX1 \fGy_tri_enable_reg[0]  ( .D(n5379), .CLK(clk), .Q(N4466) );
  DFFPOSX1 \fGy_tri_enable_reg[1]  ( .D(n5378), .CLK(clk), .Q(N4463) );
  DFFPOSX1 \fGy_tri_enable_reg[2]  ( .D(n5377), .CLK(clk), .Q(N4460) );
  DFFPOSX1 \fGy_tri_enable_reg[3]  ( .D(n5376), .CLK(clk), .Q(N4457) );
  DFFPOSX1 \fGy_tri_enable_reg[4]  ( .D(n5375), .CLK(clk), .Q(N4454) );
  DFFPOSX1 \fGy_tri_enable_reg[5]  ( .D(n5374), .CLK(clk), .Q(N4451) );
  DFFPOSX1 \fGy_tri_enable_reg[6]  ( .D(n5373), .CLK(clk), .Q(N4448) );
  DFFPOSX1 \fGy_tri_enable_reg[7]  ( .D(n5372), .CLK(clk), .Q(N4445) );
  DFFPOSX1 \fGx_tri_enable_reg[7]  ( .D(n5371), .CLK(clk), .Q(N4373) );
  DFFPOSX1 \fGx_tri_enable_reg[6]  ( .D(n5370), .CLK(clk), .Q(N4376) );
  DFFPOSX1 \fGx_tri_enable_reg[5]  ( .D(n5369), .CLK(clk), .Q(N4379) );
  DFFPOSX1 \fGx_tri_enable_reg[4]  ( .D(n5368), .CLK(clk), .Q(N4382) );
  DFFPOSX1 \fGx_tri_enable_reg[3]  ( .D(n5367), .CLK(clk), .Q(N4385) );
  DFFPOSX1 \fGx_tri_enable_reg[2]  ( .D(n5366), .CLK(clk), .Q(N4388) );
  DFFPOSX1 \fGx_tri_enable_reg[1]  ( .D(n5365), .CLK(clk), .Q(N4391) );
  DFFPOSX1 \fGx_tri_enable_reg[0]  ( .D(n5364), .CLK(clk), .Q(N4394) );
  DFFPOSX1 \dx_tri_enable_reg[0]  ( .D(n5363), .CLK(clk), .Q(N4502) );
  DFFPOSX1 \regX_reg[15][0]  ( .D(n5362), .CLK(clk), .Q(\regX[15][0] ) );
  DFFPOSX1 \regX_reg[15][1]  ( .D(n5361), .CLK(clk), .Q(\regX[15][1] ) );
  DFFPOSX1 \regX_reg[15][2]  ( .D(n5360), .CLK(clk), .Q(\regX[15][2] ) );
  DFFPOSX1 \regX_reg[15][3]  ( .D(n5359), .CLK(clk), .Q(\regX[15][3] ) );
  DFFPOSX1 \regX_reg[15][4]  ( .D(n5358), .CLK(clk), .Q(\regX[15][4] ) );
  DFFPOSX1 \regX_reg[15][5]  ( .D(n5357), .CLK(clk), .Q(\regX[15][5] ) );
  DFFPOSX1 \regX_reg[15][6]  ( .D(n5356), .CLK(clk), .Q(\regX[15][6] ) );
  DFFPOSX1 \regX_reg[15][7]  ( .D(n5355), .CLK(clk), .Q(\regX[15][7] ) );
  DFFPOSX1 \regX_reg[0][2]  ( .D(n5354), .CLK(clk), .Q(\regX[0][2] ) );
  DFFPOSX1 \regX_reg[0][3]  ( .D(n5353), .CLK(clk), .Q(\regX[0][3] ) );
  DFFPOSX1 \regX_reg[0][4]  ( .D(n5352), .CLK(clk), .Q(\regX[0][4] ) );
  DFFPOSX1 \regX_reg[0][5]  ( .D(n5351), .CLK(clk), .Q(\regX[0][5] ) );
  DFFPOSX1 \regX_reg[0][6]  ( .D(n5350), .CLK(clk), .Q(\regX[0][6] ) );
  DFFPOSX1 \regX_reg[0][7]  ( .D(n5349), .CLK(clk), .Q(\regX[0][7] ) );
  DFFPOSX1 \regX_reg[0][1]  ( .D(n5348), .CLK(clk), .Q(\regX[0][1] ) );
  DFFPOSX1 \regX_reg[0][0]  ( .D(n5347), .CLK(clk), .Q(\regX[0][0] ) );
  DFFPOSX1 \regX_reg[13][7]  ( .D(n5346), .CLK(clk), .Q(\regX[13][7] ) );
  DFFPOSX1 \regX_reg[13][6]  ( .D(n5345), .CLK(clk), .Q(\regX[13][6] ) );
  DFFPOSX1 \regX_reg[13][5]  ( .D(n5344), .CLK(clk), .Q(\regX[13][5] ) );
  DFFPOSX1 \regX_reg[13][4]  ( .D(n5343), .CLK(clk), .Q(\regX[13][4] ) );
  DFFPOSX1 \regX_reg[13][3]  ( .D(n5342), .CLK(clk), .Q(\regX[13][3] ) );
  DFFPOSX1 \regX_reg[13][2]  ( .D(n5341), .CLK(clk), .Q(\regX[13][2] ) );
  DFFPOSX1 \regX_reg[13][1]  ( .D(n5340), .CLK(clk), .Q(\regX[13][1] ) );
  DFFPOSX1 \regX_reg[13][0]  ( .D(n5339), .CLK(clk), .Q(\regX[13][0] ) );
  DFFPOSX1 \regZ_reg[12][0]  ( .D(n5338), .CLK(clk), .Q(N4081) );
  DFFPOSX1 \regZ_tri_enable_reg[12][0]  ( .D(n5337), .CLK(clk), .Q(N4082) );
  DFFPOSX1 \regZ_tri_enable_reg[12][7]  ( .D(n5336), .CLK(clk), .Q(N4061) );
  DFFPOSX1 \regZ_reg[12][7]  ( .D(n5335), .CLK(clk), .Q(N4060) );
  DFFPOSX1 \regZ_tri_enable_reg[12][6]  ( .D(n5334), .CLK(clk), .Q(N4064) );
  DFFPOSX1 \regZ_reg[12][6]  ( .D(n5333), .CLK(clk), .Q(N4063) );
  DFFPOSX1 \regZ_tri_enable_reg[12][5]  ( .D(n5332), .CLK(clk), .Q(N4067) );
  DFFPOSX1 \regZ_reg[12][5]  ( .D(n5331), .CLK(clk), .Q(N4066) );
  DFFPOSX1 \regZ_tri_enable_reg[12][4]  ( .D(n5330), .CLK(clk), .Q(N4070) );
  DFFPOSX1 \regZ_reg[12][4]  ( .D(n5329), .CLK(clk), .Q(N4069) );
  DFFPOSX1 \regZ_tri_enable_reg[12][3]  ( .D(n5328), .CLK(clk), .Q(N4073) );
  DFFPOSX1 \regZ_reg[12][3]  ( .D(n5327), .CLK(clk), .Q(N4072) );
  DFFPOSX1 \regZ_tri_enable_reg[12][2]  ( .D(n5326), .CLK(clk), .Q(N4076) );
  DFFPOSX1 \regZ_reg[12][2]  ( .D(n5325), .CLK(clk), .Q(N4075) );
  DFFPOSX1 \regZ_tri_enable_reg[12][1]  ( .D(n5324), .CLK(clk), .Q(N4079) );
  DFFPOSX1 \regZ_reg[12][1]  ( .D(n5323), .CLK(clk), .Q(N4078) );
  DFFPOSX1 \regZ_reg[0][0]  ( .D(n5322), .CLK(clk), .Q(N3793) );
  DFFPOSX1 \regZ_tri_enable_reg[0][0]  ( .D(n5321), .CLK(clk), .Q(N3794) );
  DFFPOSX1 \regZ_reg[0][1]  ( .D(n5320), .CLK(clk), .Q(N3790) );
  DFFPOSX1 \regZ_tri_enable_reg[0][1]  ( .D(n5319), .CLK(clk), .Q(N3791) );
  DFFPOSX1 \regZ_reg[0][2]  ( .D(n5318), .CLK(clk), .Q(N3787) );
  DFFPOSX1 \regZ_tri_enable_reg[0][2]  ( .D(n5317), .CLK(clk), .Q(N3788) );
  DFFPOSX1 \regZ_reg[0][3]  ( .D(n5316), .CLK(clk), .Q(N3784) );
  DFFPOSX1 \regZ_tri_enable_reg[0][3]  ( .D(n5315), .CLK(clk), .Q(N3785) );
  DFFPOSX1 \regZ_tri_enable_reg[0][7]  ( .D(n5314), .CLK(clk), .Q(N3773) );
  DFFPOSX1 \regZ_reg[0][7]  ( .D(n5313), .CLK(clk), .Q(N3772) );
  DFFPOSX1 \regZ_tri_enable_reg[0][6]  ( .D(n5312), .CLK(clk), .Q(N3776) );
  DFFPOSX1 \regZ_reg[0][6]  ( .D(n5311), .CLK(clk), .Q(N3775) );
  DFFPOSX1 \regZ_tri_enable_reg[0][5]  ( .D(n5310), .CLK(clk), .Q(N3779) );
  DFFPOSX1 \regZ_reg[0][5]  ( .D(n5309), .CLK(clk), .Q(N3778) );
  DFFPOSX1 \regZ_tri_enable_reg[0][4]  ( .D(n5308), .CLK(clk), .Q(N3782) );
  DFFPOSX1 \regZ_reg[0][4]  ( .D(n5307), .CLK(clk), .Q(N3781) );
  DFFPOSX1 \regY_reg[6][0]  ( .D(n12446), .CLK(clk), .Q(\regY[6][0] ) );
  DFFPOSX1 \regY_reg[6][1]  ( .D(n8291), .CLK(clk), .Q(\regY[6][1] ) );
  DFFPOSX1 \regY_reg[6][2]  ( .D(n12447), .CLK(clk), .Q(\regY[6][2] ) );
  DFFPOSX1 \regY_reg[6][3]  ( .D(n8289), .CLK(clk), .Q(\regY[6][3] ) );
  DFFPOSX1 \regY_reg[6][4]  ( .D(n8288), .CLK(clk), .Q(\regY[6][4] ) );
  DFFPOSX1 \regY_reg[6][5]  ( .D(n8287), .CLK(clk), .Q(\regY[6][5] ) );
  DFFPOSX1 \regY_reg[6][6]  ( .D(n15324), .CLK(clk), .Q(\regY[6][6] ) );
  DFFPOSX1 \regY_reg[6][7]  ( .D(n15323), .CLK(clk), .Q(\regY[6][7] ) );
  DFFPOSX1 \dx_reg[1]  ( .D(n8314), .CLK(clk), .Q(dx[1]) );
  DFFPOSX1 \dy_reg[1]  ( .D(n5297), .CLK(clk), .Q(dy[1]) );
  DFFPOSX1 \dx_reg[0]  ( .D(n5296), .CLK(clk), .Q(N4501) );
  DFFPOSX1 \dy_reg[0]  ( .D(n5295), .CLK(clk), .Q(N4495) );
  DFFPOSX1 \dy_tri_enable_reg[0]  ( .D(n5294), .CLK(clk), .Q(N4496) );
  DFFPOSX1 \regX_reg[6][0]  ( .D(n5293), .CLK(clk), .Q(\regX[6][0] ) );
  DFFPOSX1 \regX_reg[6][1]  ( .D(n5292), .CLK(clk), .Q(\regX[6][1] ) );
  DFFPOSX1 \regX_reg[6][2]  ( .D(n5291), .CLK(clk), .Q(\regX[6][2] ) );
  DFFPOSX1 \regX_reg[6][3]  ( .D(n5290), .CLK(clk), .Q(\regX[6][3] ) );
  DFFPOSX1 \regX_reg[6][4]  ( .D(n5289), .CLK(clk), .Q(\regX[6][4] ) );
  DFFPOSX1 \regX_reg[6][5]  ( .D(n5288), .CLK(clk), .Q(\regX[6][5] ) );
  DFFPOSX1 \regX_reg[6][6]  ( .D(n5287), .CLK(clk), .Q(\regX[6][6] ) );
  DFFPOSX1 \regX_reg[6][7]  ( .D(n5286), .CLK(clk), .Q(\regX[6][7] ) );
  DFFPOSX1 \regX_reg[1][0]  ( .D(n5285), .CLK(clk), .Q(\regX[1][0] ) );
  DFFPOSX1 \regX_reg[1][1]  ( .D(n5284), .CLK(clk), .Q(\regX[1][1] ) );
  DFFPOSX1 \regX_reg[1][2]  ( .D(n5283), .CLK(clk), .Q(\regX[1][2] ) );
  DFFPOSX1 \regX_reg[1][3]  ( .D(n5282), .CLK(clk), .Q(\regX[1][3] ) );
  DFFPOSX1 \regX_reg[1][4]  ( .D(n5281), .CLK(clk), .Q(\regX[1][4] ) );
  DFFPOSX1 \regX_reg[1][5]  ( .D(n5280), .CLK(clk), .Q(\regX[1][5] ) );
  DFFPOSX1 \regX_reg[1][6]  ( .D(n5279), .CLK(clk), .Q(\regX[1][6] ) );
  DFFPOSX1 \regX_reg[1][7]  ( .D(n5278), .CLK(clk), .Q(\regX[1][7] ) );
  DFFPOSX1 \regX_reg[2][0]  ( .D(n5277), .CLK(clk), .Q(N1375) );
  DFFPOSX1 \regX_reg[2][1]  ( .D(n5276), .CLK(clk), .Q(N1376) );
  DFFPOSX1 \regX_reg[2][2]  ( .D(n5275), .CLK(clk), .Q(N1377) );
  DFFPOSX1 \regX_reg[2][3]  ( .D(n5274), .CLK(clk), .Q(N1378) );
  DFFPOSX1 \regX_reg[2][4]  ( .D(n5273), .CLK(clk), .Q(N1379) );
  DFFPOSX1 \regX_reg[2][5]  ( .D(n5272), .CLK(clk), .Q(N1380) );
  DFFPOSX1 \regX_reg[2][6]  ( .D(n5271), .CLK(clk), .Q(N1381) );
  DFFPOSX1 \regX_reg[2][7]  ( .D(n5270), .CLK(clk), .Q(N1382) );
  DFFPOSX1 \regX_reg[3][0]  ( .D(n5269), .CLK(clk), .Q(\regX[3][0] ) );
  DFFPOSX1 \regX_reg[3][1]  ( .D(n5268), .CLK(clk), .Q(\regX[3][1] ) );
  DFFPOSX1 \regX_reg[3][2]  ( .D(n5267), .CLK(clk), .Q(\regX[3][2] ) );
  DFFPOSX1 \regX_reg[3][3]  ( .D(n5266), .CLK(clk), .Q(\regX[3][3] ) );
  DFFPOSX1 \regX_reg[3][4]  ( .D(n5265), .CLK(clk), .Q(\regX[3][4] ) );
  DFFPOSX1 \regX_reg[3][5]  ( .D(n5264), .CLK(clk), .Q(\regX[3][5] ) );
  DFFPOSX1 \regX_reg[3][6]  ( .D(n5263), .CLK(clk), .Q(\regX[3][6] ) );
  DFFPOSX1 \regX_reg[3][7]  ( .D(n5262), .CLK(clk), .Q(\regX[3][7] ) );
  DFFPOSX1 \regX_reg[4][0]  ( .D(n5261), .CLK(clk), .Q(N1433) );
  DFFPOSX1 \regX_reg[4][1]  ( .D(n5260), .CLK(clk), .Q(N1434) );
  DFFPOSX1 \regX_reg[4][2]  ( .D(n5259), .CLK(clk), .Q(N1435) );
  DFFPOSX1 \regX_reg[4][3]  ( .D(n5258), .CLK(clk), .Q(N1436) );
  DFFPOSX1 \regX_reg[4][4]  ( .D(n5257), .CLK(clk), .Q(N1437) );
  DFFPOSX1 \regX_reg[4][5]  ( .D(n5256), .CLK(clk), .Q(N1438) );
  DFFPOSX1 \regX_reg[4][6]  ( .D(n5255), .CLK(clk), .Q(N1439) );
  DFFPOSX1 \regX_reg[4][7]  ( .D(n5254), .CLK(clk), .Q(N1440) );
  DFFPOSX1 \regX_reg[5][0]  ( .D(n5253), .CLK(clk), .Q(\regX[5][0] ) );
  DFFPOSX1 \regX_reg[5][1]  ( .D(n5252), .CLK(clk), .Q(\regX[5][1] ) );
  DFFPOSX1 \regX_reg[5][2]  ( .D(n5251), .CLK(clk), .Q(\regX[5][2] ) );
  DFFPOSX1 \regX_reg[5][3]  ( .D(n5250), .CLK(clk), .Q(\regX[5][3] ) );
  DFFPOSX1 \regX_reg[5][4]  ( .D(n5249), .CLK(clk), .Q(\regX[5][4] ) );
  DFFPOSX1 \regX_reg[5][5]  ( .D(n5248), .CLK(clk), .Q(\regX[5][5] ) );
  DFFPOSX1 \regX_reg[5][6]  ( .D(n5247), .CLK(clk), .Q(\regX[5][6] ) );
  DFFPOSX1 \regX_reg[5][7]  ( .D(n5246), .CLK(clk), .Q(\regX[5][7] ) );
  DFFPOSX1 \regX_reg[7][0]  ( .D(n5245), .CLK(clk), .Q(\regX[7][0] ) );
  DFFPOSX1 \regX_reg[7][1]  ( .D(n5244), .CLK(clk), .Q(\regX[7][1] ) );
  DFFPOSX1 \regX_reg[7][2]  ( .D(n5243), .CLK(clk), .Q(\regX[7][2] ) );
  DFFPOSX1 \regX_reg[7][3]  ( .D(n5242), .CLK(clk), .Q(\regX[7][3] ) );
  DFFPOSX1 \regX_reg[7][4]  ( .D(n5241), .CLK(clk), .Q(\regX[7][4] ) );
  DFFPOSX1 \regX_reg[7][5]  ( .D(n5240), .CLK(clk), .Q(\regX[7][5] ) );
  DFFPOSX1 \regX_reg[7][6]  ( .D(n5239), .CLK(clk), .Q(\regX[7][6] ) );
  DFFPOSX1 \regX_reg[7][7]  ( .D(n5238), .CLK(clk), .Q(\regX[7][7] ) );
  DFFPOSX1 \regX_reg[8][0]  ( .D(n5237), .CLK(clk), .Q(\regX[8][0] ) );
  DFFPOSX1 \regX_reg[8][1]  ( .D(n5236), .CLK(clk), .Q(\regX[8][1] ) );
  DFFPOSX1 \regX_reg[8][2]  ( .D(n5235), .CLK(clk), .Q(\regX[8][2] ) );
  DFFPOSX1 \regX_reg[8][3]  ( .D(n5234), .CLK(clk), .Q(\regX[8][3] ) );
  DFFPOSX1 \regX_reg[8][4]  ( .D(n5233), .CLK(clk), .Q(\regX[8][4] ) );
  DFFPOSX1 \regX_reg[8][5]  ( .D(n5232), .CLK(clk), .Q(\regX[8][5] ) );
  DFFPOSX1 \regX_reg[8][6]  ( .D(n5231), .CLK(clk), .Q(\regX[8][6] ) );
  DFFPOSX1 \regX_reg[8][7]  ( .D(n5230), .CLK(clk), .Q(\regX[8][7] ) );
  DFFPOSX1 \regX_reg[9][0]  ( .D(n5229), .CLK(clk), .Q(\regX[9][0] ) );
  DFFPOSX1 \regX_reg[9][1]  ( .D(n5228), .CLK(clk), .Q(\regX[9][1] ) );
  DFFPOSX1 \regX_reg[9][2]  ( .D(n5227), .CLK(clk), .Q(\regX[9][2] ) );
  DFFPOSX1 \regX_reg[9][3]  ( .D(n5226), .CLK(clk), .Q(\regX[9][3] ) );
  DFFPOSX1 \regX_reg[9][4]  ( .D(n5225), .CLK(clk), .Q(\regX[9][4] ) );
  DFFPOSX1 \regX_reg[9][5]  ( .D(n5224), .CLK(clk), .Q(\regX[9][5] ) );
  DFFPOSX1 \regX_reg[9][6]  ( .D(n5223), .CLK(clk), .Q(\regX[9][6] ) );
  DFFPOSX1 \regX_reg[9][7]  ( .D(n5222), .CLK(clk), .Q(\regX[9][7] ) );
  DFFPOSX1 \regX_reg[16][0]  ( .D(n5221), .CLK(clk), .Q(\regX[16][0] ) );
  DFFPOSX1 \regX_reg[16][1]  ( .D(n5220), .CLK(clk), .Q(\regX[16][1] ) );
  DFFPOSX1 \regX_reg[16][2]  ( .D(n5219), .CLK(clk), .Q(\regX[16][2] ) );
  DFFPOSX1 \regX_reg[16][3]  ( .D(n5218), .CLK(clk), .Q(\regX[16][3] ) );
  DFFPOSX1 \regX_reg[16][4]  ( .D(n5217), .CLK(clk), .Q(\regX[16][4] ) );
  DFFPOSX1 \regX_reg[16][5]  ( .D(n5216), .CLK(clk), .Q(\regX[16][5] ) );
  DFFPOSX1 \regX_reg[16][6]  ( .D(n5215), .CLK(clk), .Q(\regX[16][6] ) );
  DFFPOSX1 \regX_reg[16][7]  ( .D(n5214), .CLK(clk), .Q(\regX[16][7] ) );
  DFFPOSX1 \regX_reg[17][0]  ( .D(n5213), .CLK(clk), .Q(\regX[17][0] ) );
  DFFPOSX1 \regX_reg[17][1]  ( .D(n5212), .CLK(clk), .Q(\regX[17][1] ) );
  DFFPOSX1 \regX_reg[17][2]  ( .D(n5211), .CLK(clk), .Q(\regX[17][2] ) );
  DFFPOSX1 \regX_reg[17][3]  ( .D(n5210), .CLK(clk), .Q(\regX[17][3] ) );
  DFFPOSX1 \regX_reg[17][4]  ( .D(n5209), .CLK(clk), .Q(\regX[17][4] ) );
  DFFPOSX1 \regX_reg[17][5]  ( .D(n5208), .CLK(clk), .Q(\regX[17][5] ) );
  DFFPOSX1 \regX_reg[17][6]  ( .D(n5207), .CLK(clk), .Q(\regX[17][6] ) );
  DFFPOSX1 \regX_reg[17][7]  ( .D(n5206), .CLK(clk), .Q(\regX[17][7] ) );
  DFFPOSX1 \regX_reg[24][0]  ( .D(n5205), .CLK(clk), .Q(\regX[24][0] ) );
  DFFPOSX1 \regX_reg[24][1]  ( .D(n5204), .CLK(clk), .Q(\regX[24][1] ) );
  DFFPOSX1 \regX_reg[24][2]  ( .D(n5203), .CLK(clk), .Q(\regX[24][2] ) );
  DFFPOSX1 \regX_reg[24][3]  ( .D(n5202), .CLK(clk), .Q(\regX[24][3] ) );
  DFFPOSX1 \regX_reg[24][4]  ( .D(n5201), .CLK(clk), .Q(\regX[24][4] ) );
  DFFPOSX1 \regX_reg[24][5]  ( .D(n5200), .CLK(clk), .Q(\regX[24][5] ) );
  DFFPOSX1 \regX_reg[24][6]  ( .D(n5199), .CLK(clk), .Q(\regX[24][6] ) );
  DFFPOSX1 \regX_reg[24][7]  ( .D(n5198), .CLK(clk), .Q(\regX[24][7] ) );
  DFFPOSX1 \regX_reg[14][0]  ( .D(n5197), .CLK(clk), .Q(N1735) );
  DFFPOSX1 \regX_reg[14][1]  ( .D(n5196), .CLK(clk), .Q(N1736) );
  DFFPOSX1 \regX_reg[14][2]  ( .D(n5195), .CLK(clk), .Q(N1737) );
  DFFPOSX1 \regX_reg[14][3]  ( .D(n5194), .CLK(clk), .Q(N1738) );
  DFFPOSX1 \regX_reg[14][4]  ( .D(n5193), .CLK(clk), .Q(N1739) );
  DFFPOSX1 \regX_reg[14][5]  ( .D(n5192), .CLK(clk), .Q(N1740) );
  DFFPOSX1 \regX_reg[14][6]  ( .D(n5191), .CLK(clk), .Q(N1741) );
  DFFPOSX1 \regX_reg[14][7]  ( .D(n5190), .CLK(clk), .Q(N1742) );
  DFFPOSX1 \regX_reg[22][0]  ( .D(n5189), .CLK(clk), .Q(\regX[22][0] ) );
  DFFPOSX1 \regX_reg[22][1]  ( .D(n5188), .CLK(clk), .Q(\regX[22][1] ) );
  DFFPOSX1 \regX_reg[22][2]  ( .D(n5187), .CLK(clk), .Q(\regX[22][2] ) );
  DFFPOSX1 \regX_reg[22][3]  ( .D(n5186), .CLK(clk), .Q(\regX[22][3] ) );
  DFFPOSX1 \regX_reg[22][4]  ( .D(n5185), .CLK(clk), .Q(\regX[22][4] ) );
  DFFPOSX1 \regX_reg[22][5]  ( .D(n5184), .CLK(clk), .Q(\regX[22][5] ) );
  DFFPOSX1 \regX_reg[22][6]  ( .D(n5183), .CLK(clk), .Q(\regX[22][6] ) );
  DFFPOSX1 \regX_reg[22][7]  ( .D(n5182), .CLK(clk), .Q(\regX[22][7] ) );
  DFFPOSX1 \regX_reg[23][0]  ( .D(n5181), .CLK(clk), .Q(\regX[23][0] ) );
  DFFPOSX1 \regX_reg[23][1]  ( .D(n5180), .CLK(clk), .Q(\regX[23][1] ) );
  DFFPOSX1 \regX_reg[23][2]  ( .D(n5179), .CLK(clk), .Q(\regX[23][2] ) );
  DFFPOSX1 \regX_reg[23][3]  ( .D(n5178), .CLK(clk), .Q(\regX[23][3] ) );
  DFFPOSX1 \regX_reg[23][4]  ( .D(n5177), .CLK(clk), .Q(\regX[23][4] ) );
  DFFPOSX1 \regX_reg[23][5]  ( .D(n5176), .CLK(clk), .Q(\regX[23][5] ) );
  DFFPOSX1 \regX_reg[23][6]  ( .D(n5175), .CLK(clk), .Q(\regX[23][6] ) );
  DFFPOSX1 \regX_reg[23][7]  ( .D(n5174), .CLK(clk), .Q(\regX[23][7] ) );
  DFFPOSX1 \regX_reg[12][0]  ( .D(n5173), .CLK(clk), .Q(N1677) );
  DFFPOSX1 \regX_reg[12][1]  ( .D(n5172), .CLK(clk), .Q(N1678) );
  DFFPOSX1 \regX_reg[12][2]  ( .D(n5171), .CLK(clk), .Q(N1679) );
  DFFPOSX1 \regX_reg[12][3]  ( .D(n5170), .CLK(clk), .Q(N1680) );
  DFFPOSX1 \regX_reg[12][4]  ( .D(n5169), .CLK(clk), .Q(N1681) );
  DFFPOSX1 \regX_reg[12][5]  ( .D(n5168), .CLK(clk), .Q(N1682) );
  DFFPOSX1 \regX_reg[12][6]  ( .D(n5167), .CLK(clk), .Q(N1683) );
  DFFPOSX1 \regX_reg[12][7]  ( .D(n5166), .CLK(clk), .Q(N1684) );
  DFFPOSX1 \regX_reg[20][0]  ( .D(n5165), .CLK(clk), .Q(\regX[20][0] ) );
  DFFPOSX1 \regX_reg[20][1]  ( .D(n5164), .CLK(clk), .Q(\regX[20][1] ) );
  DFFPOSX1 \regX_reg[20][2]  ( .D(n5163), .CLK(clk), .Q(\regX[20][2] ) );
  DFFPOSX1 \regX_reg[20][3]  ( .D(n5162), .CLK(clk), .Q(\regX[20][3] ) );
  DFFPOSX1 \regX_reg[20][4]  ( .D(n5161), .CLK(clk), .Q(\regX[20][4] ) );
  DFFPOSX1 \regX_reg[20][5]  ( .D(n5160), .CLK(clk), .Q(\regX[20][5] ) );
  DFFPOSX1 \regX_reg[20][6]  ( .D(n5159), .CLK(clk), .Q(\regX[20][6] ) );
  DFFPOSX1 \regX_reg[20][7]  ( .D(n5158), .CLK(clk), .Q(\regX[20][7] ) );
  DFFPOSX1 \regX_reg[21][0]  ( .D(n5157), .CLK(clk), .Q(\regX[21][0] ) );
  DFFPOSX1 \regX_reg[21][1]  ( .D(n5156), .CLK(clk), .Q(\regX[21][1] ) );
  DFFPOSX1 \regX_reg[21][2]  ( .D(n5155), .CLK(clk), .Q(\regX[21][2] ) );
  DFFPOSX1 \regX_reg[21][3]  ( .D(n5154), .CLK(clk), .Q(\regX[21][3] ) );
  DFFPOSX1 \regX_reg[21][4]  ( .D(n5153), .CLK(clk), .Q(\regX[21][4] ) );
  DFFPOSX1 \regX_reg[21][5]  ( .D(n5152), .CLK(clk), .Q(\regX[21][5] ) );
  DFFPOSX1 \regX_reg[21][6]  ( .D(n5151), .CLK(clk), .Q(\regX[21][6] ) );
  DFFPOSX1 \regX_reg[21][7]  ( .D(n5150), .CLK(clk), .Q(\regX[21][7] ) );
  DFFPOSX1 \regX_reg[10][0]  ( .D(n5149), .CLK(clk), .Q(N1615) );
  DFFPOSX1 \regX_reg[10][1]  ( .D(n5148), .CLK(clk), .Q(N1616) );
  DFFPOSX1 \regX_reg[10][2]  ( .D(n5147), .CLK(clk), .Q(N1617) );
  DFFPOSX1 \regX_reg[10][3]  ( .D(n5146), .CLK(clk), .Q(N1618) );
  DFFPOSX1 \regX_reg[10][4]  ( .D(n5145), .CLK(clk), .Q(N1619) );
  DFFPOSX1 \regX_reg[10][5]  ( .D(n5144), .CLK(clk), .Q(N1620) );
  DFFPOSX1 \regX_reg[10][6]  ( .D(n5143), .CLK(clk), .Q(N1621) );
  DFFPOSX1 \regX_reg[10][7]  ( .D(n5142), .CLK(clk), .Q(N1622) );
  DFFPOSX1 \regX_reg[11][0]  ( .D(n5141), .CLK(clk), .Q(\regX[11][0] ) );
  DFFPOSX1 \regX_reg[11][1]  ( .D(n5140), .CLK(clk), .Q(\regX[11][1] ) );
  DFFPOSX1 \regX_reg[11][2]  ( .D(n5139), .CLK(clk), .Q(\regX[11][2] ) );
  DFFPOSX1 \regX_reg[11][3]  ( .D(n5138), .CLK(clk), .Q(\regX[11][3] ) );
  DFFPOSX1 \regX_reg[11][4]  ( .D(n5137), .CLK(clk), .Q(\regX[11][4] ) );
  DFFPOSX1 \regX_reg[11][5]  ( .D(n5136), .CLK(clk), .Q(\regX[11][5] ) );
  DFFPOSX1 \regX_reg[11][6]  ( .D(n5135), .CLK(clk), .Q(\regX[11][6] ) );
  DFFPOSX1 \regX_reg[11][7]  ( .D(n5134), .CLK(clk), .Q(\regX[11][7] ) );
  DFFPOSX1 \Gy_reg[0]  ( .D(n5133), .CLK(clk), .Q(Gy[0]) );
  DFFPOSX1 \Gy_reg[1]  ( .D(n5132), .CLK(clk), .Q(Gy[1]) );
  DFFPOSX1 \Gy_reg[2]  ( .D(n5131), .CLK(clk), .Q(Gy[2]) );
  DFFPOSX1 \Gy_reg[3]  ( .D(n5130), .CLK(clk), .Q(Gy[3]) );
  DFFPOSX1 \Gy_reg[4]  ( .D(n5129), .CLK(clk), .Q(Gy[4]) );
  DFFPOSX1 \Gy_reg[5]  ( .D(n5128), .CLK(clk), .Q(Gy[5]) );
  DFFPOSX1 \Gy_reg[6]  ( .D(n5127), .CLK(clk), .Q(Gy[6]) );
  DFFPOSX1 \Gy_reg[7]  ( .D(n5126), .CLK(clk), .Q(Gy[7]) );
  DFFPOSX1 \Gy_reg[8]  ( .D(n5125), .CLK(clk), .Q(Gy[8]) );
  DFFPOSX1 \Gy_reg[9]  ( .D(n5124), .CLK(clk), .Q(Gy[9]) );
  DFFPOSX1 \Gy_reg[10]  ( .D(n5123), .CLK(clk), .Q(Gy[10]) );
  DFFPOSX1 \Gy_reg[11]  ( .D(n5122), .CLK(clk), .Q(Gy[11]) );
  DFFPOSX1 \Gy_reg[12]  ( .D(n5121), .CLK(clk), .Q(Gy[12]) );
  DFFPOSX1 \Gy_reg[13]  ( .D(n5120), .CLK(clk), .Q(Gy[13]) );
  DFFPOSX1 \Gy_reg[14]  ( .D(n5119), .CLK(clk), .Q(Gy[14]) );
  DFFPOSX1 \Gy_reg[15]  ( .D(n5118), .CLK(clk), .Q(Gy[15]) );
  DFFPOSX1 \Gy_reg[16]  ( .D(n5117), .CLK(clk), .Q(Gy[16]) );
  DFFPOSX1 \Gy_reg[17]  ( .D(n5116), .CLK(clk), .Q(Gy[17]) );
  DFFPOSX1 \Gy_reg[18]  ( .D(n5115), .CLK(clk), .Q(Gy[18]) );
  DFFPOSX1 \Gy_reg[19]  ( .D(n5114), .CLK(clk), .Q(Gy[19]) );
  DFFPOSX1 \Gy_reg[20]  ( .D(n5113), .CLK(clk), .Q(Gy[20]) );
  DFFPOSX1 \Gy_reg[21]  ( .D(n5112), .CLK(clk), .Q(Gy[21]) );
  DFFPOSX1 \Gy_reg[22]  ( .D(n5111), .CLK(clk), .Q(Gy[22]) );
  DFFPOSX1 \Gy_reg[23]  ( .D(n5110), .CLK(clk), .Q(Gy[23]) );
  DFFPOSX1 \Gy_reg[24]  ( .D(n5109), .CLK(clk), .Q(Gy[24]) );
  DFFPOSX1 \Gy_reg[25]  ( .D(n5108), .CLK(clk), .Q(Gy[25]) );
  DFFPOSX1 \Gy_reg[26]  ( .D(n5107), .CLK(clk), .Q(Gy[26]) );
  DFFPOSX1 \Gy_reg[27]  ( .D(n5106), .CLK(clk), .Q(Gy[27]) );
  DFFPOSX1 \Gy_reg[28]  ( .D(n5105), .CLK(clk), .Q(Gy[28]) );
  DFFPOSX1 \Gy_reg[29]  ( .D(n5104), .CLK(clk), .Q(Gy[29]) );
  DFFPOSX1 \Gy_reg[30]  ( .D(n5103), .CLK(clk), .Q(Gy[30]) );
  DFFPOSX1 \Gy_reg[31]  ( .D(n5102), .CLK(clk), .Q(Gy[31]) );
  DFFPOSX1 \Out_gradient_tri_enable_reg[0]  ( .D(n5101), .CLK(clk), .Q(N4418)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[1]  ( .D(n5100), .CLK(clk), .Q(N4415)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[2]  ( .D(n5099), .CLK(clk), .Q(N4412)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[3]  ( .D(n5098), .CLK(clk), .Q(N4409)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[4]  ( .D(n5097), .CLK(clk), .Q(N4406)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[5]  ( .D(n5096), .CLK(clk), .Q(N4403)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[6]  ( .D(n5095), .CLK(clk), .Q(N4400)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[7]  ( .D(n5094), .CLK(clk), .Q(N4397)
         );
  DFFPOSX1 \fGx_reg[8]  ( .D(n5093), .CLK(clk), .Q(fGx[8]) );
  DFFPOSX1 \fGy_reg[0]  ( .D(n5092), .CLK(clk), .Q(N4465) );
  DFFPOSX1 \fGy_reg[1]  ( .D(n5091), .CLK(clk), .Q(N4462) );
  DFFPOSX1 \fGy_reg[2]  ( .D(n5090), .CLK(clk), .Q(N4459) );
  DFFPOSX1 \fGy_reg[3]  ( .D(n5089), .CLK(clk), .Q(N4456) );
  DFFPOSX1 \fGy_reg[4]  ( .D(n5088), .CLK(clk), .Q(N4453) );
  DFFPOSX1 \fGy_reg[5]  ( .D(n5087), .CLK(clk), .Q(N4450) );
  DFFPOSX1 \fGy_reg[6]  ( .D(n5086), .CLK(clk), .Q(N4447) );
  DFFPOSX1 \fGy_reg[7]  ( .D(n5085), .CLK(clk), .Q(N4444) );
  DFFPOSX1 \fGy_reg[8]  ( .D(n5084), .CLK(clk), .Q(fGy[8]) );
  DFFPOSX1 \fGy_reg[9]  ( .D(n5083), .CLK(clk), .Q(fGy[9]) );
  DFFPOSX1 \fGy_reg[10]  ( .D(n5082), .CLK(clk), .Q(fGy[10]) );
  DFFPOSX1 \fGy_reg[11]  ( .D(n5081), .CLK(clk), .Q(fGy[11]) );
  DFFPOSX1 \fGy_reg[12]  ( .D(n5080), .CLK(clk), .Q(fGy[12]) );
  DFFPOSX1 \fGy_reg[13]  ( .D(n5079), .CLK(clk), .Q(fGy[13]) );
  DFFPOSX1 \fGy_reg[14]  ( .D(n5078), .CLK(clk), .Q(fGy[14]) );
  DFFPOSX1 \fGy_reg[15]  ( .D(n5077), .CLK(clk), .Q(fGy[15]) );
  DFFPOSX1 \fGy_reg[16]  ( .D(n5076), .CLK(clk), .Q(fGy[16]) );
  DFFPOSX1 \fGy_reg[17]  ( .D(n5075), .CLK(clk), .Q(fGy[17]) );
  DFFPOSX1 \fGy_reg[18]  ( .D(n5074), .CLK(clk), .Q(fGy[18]) );
  DFFPOSX1 \fGy_reg[19]  ( .D(n5073), .CLK(clk), .Q(fGy[19]) );
  DFFPOSX1 \fGy_reg[20]  ( .D(n5072), .CLK(clk), .Q(fGy[20]) );
  DFFPOSX1 \fGy_reg[21]  ( .D(n5071), .CLK(clk), .Q(fGy[21]) );
  DFFPOSX1 \fGy_reg[22]  ( .D(n5070), .CLK(clk), .Q(fGy[22]) );
  DFFPOSX1 \fGy_reg[23]  ( .D(n5069), .CLK(clk), .Q(fGy[23]) );
  DFFPOSX1 \fGy_reg[24]  ( .D(n5068), .CLK(clk), .Q(fGy[24]) );
  DFFPOSX1 \fGy_reg[25]  ( .D(n5067), .CLK(clk), .Q(fGy[25]) );
  DFFPOSX1 \fGy_reg[26]  ( .D(n5066), .CLK(clk), .Q(fGy[26]) );
  DFFPOSX1 \fGy_reg[27]  ( .D(n5065), .CLK(clk), .Q(fGy[27]) );
  DFFPOSX1 \fGy_reg[28]  ( .D(n5064), .CLK(clk), .Q(fGy[28]) );
  DFFPOSX1 \fGy_reg[29]  ( .D(n5063), .CLK(clk), .Q(fGy[29]) );
  DFFPOSX1 \fGy_reg[30]  ( .D(n5062), .CLK(clk), .Q(fGy[30]) );
  DFFPOSX1 \fGy_reg[31]  ( .D(n5061), .CLK(clk), .Q(fGy[31]) );
  DFFPOSX1 \Gx_reg[0]  ( .D(n5060), .CLK(clk), .Q(Gx[0]) );
  DFFPOSX1 \fGx_reg[0]  ( .D(n5059), .CLK(clk), .Q(N4393) );
  DFFPOSX1 \Gx_reg[1]  ( .D(n5058), .CLK(clk), .Q(Gx[1]) );
  DFFPOSX1 \fGx_reg[1]  ( .D(n5057), .CLK(clk), .Q(N4390) );
  DFFPOSX1 \Gx_reg[2]  ( .D(n5056), .CLK(clk), .Q(Gx[2]) );
  DFFPOSX1 \fGx_reg[2]  ( .D(n5055), .CLK(clk), .Q(N4387) );
  DFFPOSX1 \Gx_reg[3]  ( .D(n5054), .CLK(clk), .Q(Gx[3]) );
  DFFPOSX1 \fGx_reg[3]  ( .D(n5053), .CLK(clk), .Q(N4384) );
  DFFPOSX1 \Gx_reg[4]  ( .D(n5052), .CLK(clk), .Q(Gx[4]) );
  DFFPOSX1 \fGx_reg[4]  ( .D(n5051), .CLK(clk), .Q(N4381) );
  DFFPOSX1 \Gx_reg[5]  ( .D(n5050), .CLK(clk), .Q(Gx[5]) );
  DFFPOSX1 \fGx_reg[5]  ( .D(n5049), .CLK(clk), .Q(N4378) );
  DFFPOSX1 \Gx_reg[6]  ( .D(n5048), .CLK(clk), .Q(Gx[6]) );
  DFFPOSX1 \fGx_reg[6]  ( .D(n5047), .CLK(clk), .Q(N4375) );
  DFFPOSX1 \Gx_reg[7]  ( .D(n5046), .CLK(clk), .Q(Gx[7]) );
  DFFPOSX1 \fGx_reg[7]  ( .D(n5045), .CLK(clk), .Q(N4372) );
  DFFPOSX1 \Gx_reg[8]  ( .D(n5044), .CLK(clk), .Q(Gx[8]) );
  DFFPOSX1 \Gx_reg[9]  ( .D(n5043), .CLK(clk), .Q(Gx[9]) );
  DFFPOSX1 \fGx_reg[9]  ( .D(n5042), .CLK(clk), .Q(fGx[9]) );
  DFFPOSX1 \Gx_reg[10]  ( .D(n5041), .CLK(clk), .Q(Gx[10]) );
  DFFPOSX1 \Out_gradient_reg[0]  ( .D(n5040), .CLK(clk), .Q(N4417) );
  DFFPOSX1 \Out_gradient_reg[1]  ( .D(n5039), .CLK(clk), .Q(N4414) );
  DFFPOSX1 \Out_gradient_reg[2]  ( .D(n5038), .CLK(clk), .Q(N4411) );
  DFFPOSX1 \Out_gradient_reg[3]  ( .D(n5037), .CLK(clk), .Q(N4408) );
  DFFPOSX1 \Out_gradient_reg[4]  ( .D(n5036), .CLK(clk), .Q(N4405) );
  DFFPOSX1 \Out_gradient_reg[5]  ( .D(n5035), .CLK(clk), .Q(N4402) );
  DFFPOSX1 \Out_gradient_reg[6]  ( .D(n5034), .CLK(clk), .Q(N4399) );
  DFFPOSX1 \Out_gradient_reg[7]  ( .D(n5033), .CLK(clk), .Q(N4396) );
  DFFPOSX1 \fGx_reg[10]  ( .D(n5032), .CLK(clk), .Q(fGx[10]) );
  DFFPOSX1 \Gx_reg[11]  ( .D(n5031), .CLK(clk), .Q(Gx[11]) );
  DFFPOSX1 \fGx_reg[11]  ( .D(n5030), .CLK(clk), .Q(fGx[11]) );
  DFFPOSX1 \Gx_reg[12]  ( .D(n5029), .CLK(clk), .Q(Gx[12]) );
  DFFPOSX1 \fGx_reg[12]  ( .D(n5028), .CLK(clk), .Q(fGx[12]) );
  DFFPOSX1 \Gx_reg[13]  ( .D(n5027), .CLK(clk), .Q(Gx[13]) );
  DFFPOSX1 \fGx_reg[13]  ( .D(n5026), .CLK(clk), .Q(fGx[13]) );
  DFFPOSX1 \Gx_reg[14]  ( .D(n5025), .CLK(clk), .Q(Gx[14]) );
  DFFPOSX1 \fGx_reg[14]  ( .D(n5024), .CLK(clk), .Q(fGx[14]) );
  DFFPOSX1 \Gx_reg[15]  ( .D(n5023), .CLK(clk), .Q(Gx[15]) );
  DFFPOSX1 \fGx_reg[15]  ( .D(n5022), .CLK(clk), .Q(fGx[15]) );
  DFFPOSX1 \Gx_reg[16]  ( .D(n5021), .CLK(clk), .Q(Gx[16]) );
  DFFPOSX1 \fGx_reg[16]  ( .D(n5020), .CLK(clk), .Q(fGx[16]) );
  DFFPOSX1 \Gx_reg[17]  ( .D(n5019), .CLK(clk), .Q(Gx[17]) );
  DFFPOSX1 \fGx_reg[17]  ( .D(n5018), .CLK(clk), .Q(fGx[17]) );
  DFFPOSX1 \Gx_reg[18]  ( .D(n5017), .CLK(clk), .Q(Gx[18]) );
  DFFPOSX1 \fGx_reg[18]  ( .D(n5016), .CLK(clk), .Q(fGx[18]) );
  DFFPOSX1 \Gx_reg[19]  ( .D(n5015), .CLK(clk), .Q(Gx[19]) );
  DFFPOSX1 \fGx_reg[19]  ( .D(n5014), .CLK(clk), .Q(fGx[19]) );
  DFFPOSX1 \Gx_reg[20]  ( .D(n5013), .CLK(clk), .Q(Gx[20]) );
  DFFPOSX1 \fGx_reg[20]  ( .D(n5012), .CLK(clk), .Q(fGx[20]) );
  DFFPOSX1 \Gx_reg[21]  ( .D(n5011), .CLK(clk), .Q(Gx[21]) );
  DFFPOSX1 \fGx_reg[21]  ( .D(n5010), .CLK(clk), .Q(fGx[21]) );
  DFFPOSX1 \Gx_reg[22]  ( .D(n5009), .CLK(clk), .Q(Gx[22]) );
  DFFPOSX1 \fGx_reg[22]  ( .D(n5008), .CLK(clk), .Q(fGx[22]) );
  DFFPOSX1 \Gx_reg[23]  ( .D(n5007), .CLK(clk), .Q(Gx[23]) );
  DFFPOSX1 \fGx_reg[23]  ( .D(n5006), .CLK(clk), .Q(fGx[23]) );
  DFFPOSX1 \Gx_reg[24]  ( .D(n5005), .CLK(clk), .Q(Gx[24]) );
  DFFPOSX1 \fGx_reg[24]  ( .D(n5004), .CLK(clk), .Q(fGx[24]) );
  DFFPOSX1 \Gx_reg[25]  ( .D(n5003), .CLK(clk), .Q(Gx[25]) );
  DFFPOSX1 \fGx_reg[25]  ( .D(n5002), .CLK(clk), .Q(fGx[25]) );
  DFFPOSX1 \Gx_reg[26]  ( .D(n5001), .CLK(clk), .Q(Gx[26]) );
  DFFPOSX1 \fGx_reg[26]  ( .D(n5000), .CLK(clk), .Q(fGx[26]) );
  DFFPOSX1 \Gx_reg[27]  ( .D(n4999), .CLK(clk), .Q(Gx[27]) );
  DFFPOSX1 \fGx_reg[27]  ( .D(n4998), .CLK(clk), .Q(fGx[27]) );
  DFFPOSX1 \Gx_reg[28]  ( .D(n4997), .CLK(clk), .Q(Gx[28]) );
  DFFPOSX1 \fGx_reg[28]  ( .D(n4996), .CLK(clk), .Q(fGx[28]) );
  DFFPOSX1 \Gx_reg[29]  ( .D(n4995), .CLK(clk), .Q(Gx[29]) );
  DFFPOSX1 \fGx_reg[29]  ( .D(n4994), .CLK(clk), .Q(fGx[29]) );
  DFFPOSX1 \Gx_reg[30]  ( .D(n4993), .CLK(clk), .Q(Gx[30]) );
  DFFPOSX1 \fGx_reg[30]  ( .D(n4992), .CLK(clk), .Q(fGx[30]) );
  DFFPOSX1 \Gx_reg[31]  ( .D(n4991), .CLK(clk), .Q(Gx[31]) );
  DFFPOSX1 \fGx_reg[31]  ( .D(n4990), .CLK(clk), .Q(fGx[31]) );
  DFFPOSX1 \regX_reg[18][0]  ( .D(n4989), .CLK(clk), .Q(\regX[18][0] ) );
  DFFPOSX1 \regX_reg[18][1]  ( .D(n4988), .CLK(clk), .Q(\regX[18][1] ) );
  DFFPOSX1 \regX_reg[18][2]  ( .D(n4987), .CLK(clk), .Q(\regX[18][2] ) );
  DFFPOSX1 \regX_reg[18][3]  ( .D(n4986), .CLK(clk), .Q(\regX[18][3] ) );
  DFFPOSX1 \regX_reg[18][4]  ( .D(n4985), .CLK(clk), .Q(\regX[18][4] ) );
  DFFPOSX1 \regX_reg[18][5]  ( .D(n4984), .CLK(clk), .Q(\regX[18][5] ) );
  DFFPOSX1 \regX_reg[18][6]  ( .D(n4983), .CLK(clk), .Q(\regX[18][6] ) );
  DFFPOSX1 \regX_reg[18][7]  ( .D(n4982), .CLK(clk), .Q(\regX[18][7] ) );
  DFFPOSX1 \regX_reg[19][0]  ( .D(n4981), .CLK(clk), .Q(\regX[19][0] ) );
  DFFPOSX1 \regX_reg[19][1]  ( .D(n4980), .CLK(clk), .Q(\regX[19][1] ) );
  DFFPOSX1 \regX_reg[19][2]  ( .D(n4979), .CLK(clk), .Q(\regX[19][2] ) );
  DFFPOSX1 \regX_reg[19][3]  ( .D(n4978), .CLK(clk), .Q(\regX[19][3] ) );
  DFFPOSX1 \regX_reg[19][4]  ( .D(n4977), .CLK(clk), .Q(\regX[19][4] ) );
  DFFPOSX1 \regX_reg[19][5]  ( .D(n4976), .CLK(clk), .Q(\regX[19][5] ) );
  DFFPOSX1 \regX_reg[19][6]  ( .D(n4975), .CLK(clk), .Q(\regX[19][6] ) );
  DFFPOSX1 \regX_reg[19][7]  ( .D(n4974), .CLK(clk), .Q(\regX[19][7] ) );
  DFFPOSX1 \Out_direction_reg[0]  ( .D(n4973), .CLK(clk), .Q(N4441) );
  DFFPOSX1 \Out_direction_tri_enable_reg[0]  ( .D(n4972), .CLK(clk), .Q(N4442)
         );
  DFFPOSX1 \Out_direction_reg[1]  ( .D(n4971), .CLK(clk), .Q(N4438) );
  DFFPOSX1 \Out_direction_tri_enable_reg[1]  ( .D(n4970), .CLK(clk), .Q(N4439)
         );
  DFFPOSX1 \Out_direction_reg[2]  ( .D(n4969), .CLK(clk), .Q(N4435) );
  DFFPOSX1 \Out_direction_tri_enable_reg[2]  ( .D(n4968), .CLK(clk), .Q(N4436)
         );
  DFFPOSX1 \Out_direction_reg[3]  ( .D(n12448), .CLK(clk), .Q(N4432) );
  DFFPOSX1 \Out_direction_tri_enable_reg[3]  ( .D(n4966), .CLK(clk), .Q(N4433)
         );
  DFFPOSX1 \Out_direction_reg[4]  ( .D(n4965), .CLK(clk), .Q(N4429) );
  DFFPOSX1 \Out_direction_tri_enable_reg[4]  ( .D(n4964), .CLK(clk), .Q(N4430)
         );
  DFFPOSX1 \Out_direction_reg[5]  ( .D(n4963), .CLK(clk), .Q(N4426) );
  DFFPOSX1 \Out_direction_tri_enable_reg[5]  ( .D(n4962), .CLK(clk), .Q(N4427)
         );
  DFFPOSX1 \Out_direction_reg[6]  ( .D(n4961), .CLK(clk), .Q(N4423) );
  DFFPOSX1 \Out_direction_tri_enable_reg[6]  ( .D(n4960), .CLK(clk), .Q(N4424)
         );
  DFFPOSX1 \Out_direction_reg[7]  ( .D(n4959), .CLK(clk), .Q(N4420) );
  DFFPOSX1 \Out_direction_tri_enable_reg[7]  ( .D(n4958), .CLK(clk), .Q(N4421)
         );
  DFFPOSX1 \regZ_reg[3][0]  ( .D(n4957), .CLK(clk), .Q(N3865) );
  DFFPOSX1 \regZ_tri_enable_reg[3][0]  ( .D(n4956), .CLK(clk), .Q(N3866) );
  DFFPOSX1 \regZ_reg[3][1]  ( .D(n4955), .CLK(clk), .Q(N3862) );
  DFFPOSX1 \regZ_tri_enable_reg[3][1]  ( .D(n4954), .CLK(clk), .Q(N3863) );
  DFFPOSX1 \regZ_reg[3][2]  ( .D(n4953), .CLK(clk), .Q(N3859) );
  DFFPOSX1 \regZ_tri_enable_reg[3][2]  ( .D(n4952), .CLK(clk), .Q(N3860) );
  DFFPOSX1 \regZ_reg[3][3]  ( .D(n4951), .CLK(clk), .Q(N3856) );
  DFFPOSX1 \regZ_tri_enable_reg[3][3]  ( .D(n4950), .CLK(clk), .Q(N3857) );
  DFFPOSX1 \regZ_reg[3][4]  ( .D(n4949), .CLK(clk), .Q(N3853) );
  DFFPOSX1 \regZ_tri_enable_reg[3][4]  ( .D(n4948), .CLK(clk), .Q(N3854) );
  DFFPOSX1 \regZ_reg[3][5]  ( .D(n4947), .CLK(clk), .Q(N3850) );
  DFFPOSX1 \regZ_tri_enable_reg[3][5]  ( .D(n4946), .CLK(clk), .Q(N3851) );
  DFFPOSX1 \regZ_reg[3][6]  ( .D(n4945), .CLK(clk), .Q(N3847) );
  DFFPOSX1 \regZ_tri_enable_reg[3][6]  ( .D(n4944), .CLK(clk), .Q(N3848) );
  DFFPOSX1 \regZ_reg[3][7]  ( .D(n4943), .CLK(clk), .Q(N3844) );
  DFFPOSX1 \regZ_tri_enable_reg[3][7]  ( .D(n4942), .CLK(clk), .Q(N3845) );
  DFFPOSX1 \regZ_reg[4][0]  ( .D(n4941), .CLK(clk), .Q(N3889) );
  DFFPOSX1 \regZ_tri_enable_reg[4][0]  ( .D(n4940), .CLK(clk), .Q(N3890) );
  DFFPOSX1 \regZ_reg[4][1]  ( .D(n4939), .CLK(clk), .Q(N3886) );
  DFFPOSX1 \regZ_tri_enable_reg[4][1]  ( .D(n4938), .CLK(clk), .Q(N3887) );
  DFFPOSX1 \regZ_reg[4][2]  ( .D(n4937), .CLK(clk), .Q(N3883) );
  DFFPOSX1 \regZ_tri_enable_reg[4][2]  ( .D(n4936), .CLK(clk), .Q(N3884) );
  DFFPOSX1 \regZ_reg[4][3]  ( .D(n4935), .CLK(clk), .Q(N3880) );
  DFFPOSX1 \regZ_tri_enable_reg[4][3]  ( .D(n4934), .CLK(clk), .Q(N3881) );
  DFFPOSX1 \regZ_reg[4][4]  ( .D(n4933), .CLK(clk), .Q(N3877) );
  DFFPOSX1 \regZ_tri_enable_reg[4][4]  ( .D(n4932), .CLK(clk), .Q(N3878) );
  DFFPOSX1 \regZ_reg[4][5]  ( .D(n4931), .CLK(clk), .Q(N3874) );
  DFFPOSX1 \regZ_tri_enable_reg[4][5]  ( .D(n4930), .CLK(clk), .Q(N3875) );
  DFFPOSX1 \regZ_reg[4][6]  ( .D(n4929), .CLK(clk), .Q(N3871) );
  DFFPOSX1 \regZ_tri_enable_reg[4][6]  ( .D(n4928), .CLK(clk), .Q(N3872) );
  DFFPOSX1 \regZ_reg[4][7]  ( .D(n4927), .CLK(clk), .Q(N3868) );
  DFFPOSX1 \regZ_tri_enable_reg[4][7]  ( .D(n4926), .CLK(clk), .Q(N3869) );
  DFFPOSX1 \regZ_reg[5][0]  ( .D(n4925), .CLK(clk), .Q(N3913) );
  DFFPOSX1 \regZ_tri_enable_reg[5][0]  ( .D(n4924), .CLK(clk), .Q(N3914) );
  DFFPOSX1 \regZ_reg[5][1]  ( .D(n4923), .CLK(clk), .Q(N3910) );
  DFFPOSX1 \regZ_tri_enable_reg[5][1]  ( .D(n4922), .CLK(clk), .Q(N3911) );
  DFFPOSX1 \regZ_reg[5][2]  ( .D(n4921), .CLK(clk), .Q(N3907) );
  DFFPOSX1 \regZ_tri_enable_reg[5][2]  ( .D(n4920), .CLK(clk), .Q(N3908) );
  DFFPOSX1 \regZ_reg[5][3]  ( .D(n4919), .CLK(clk), .Q(N3904) );
  DFFPOSX1 \regZ_tri_enable_reg[5][3]  ( .D(n4918), .CLK(clk), .Q(N3905) );
  DFFPOSX1 \regZ_reg[5][4]  ( .D(n4917), .CLK(clk), .Q(N3901) );
  DFFPOSX1 \regZ_tri_enable_reg[5][4]  ( .D(n4916), .CLK(clk), .Q(N3902) );
  DFFPOSX1 \regZ_reg[5][5]  ( .D(n4915), .CLK(clk), .Q(N3898) );
  DFFPOSX1 \regZ_tri_enable_reg[5][5]  ( .D(n4914), .CLK(clk), .Q(N3899) );
  DFFPOSX1 \regZ_reg[5][6]  ( .D(n4913), .CLK(clk), .Q(N3895) );
  DFFPOSX1 \regZ_tri_enable_reg[5][6]  ( .D(n4912), .CLK(clk), .Q(N3896) );
  DFFPOSX1 \regZ_reg[5][7]  ( .D(n4911), .CLK(clk), .Q(N3892) );
  DFFPOSX1 \regZ_tri_enable_reg[5][7]  ( .D(n4910), .CLK(clk), .Q(N3893) );
  DFFPOSX1 \regZ_reg[6][0]  ( .D(n4909), .CLK(clk), .Q(N3937) );
  DFFPOSX1 \regZ_tri_enable_reg[6][0]  ( .D(n4908), .CLK(clk), .Q(N3938) );
  DFFPOSX1 \regZ_reg[6][1]  ( .D(n4907), .CLK(clk), .Q(N3934) );
  DFFPOSX1 \regZ_tri_enable_reg[6][1]  ( .D(n4906), .CLK(clk), .Q(N3935) );
  DFFPOSX1 \regZ_reg[6][2]  ( .D(n4905), .CLK(clk), .Q(N3931) );
  DFFPOSX1 \regZ_tri_enable_reg[6][2]  ( .D(n4904), .CLK(clk), .Q(N3932) );
  DFFPOSX1 \regZ_reg[6][3]  ( .D(n4903), .CLK(clk), .Q(N3928) );
  DFFPOSX1 \regZ_tri_enable_reg[6][3]  ( .D(n4902), .CLK(clk), .Q(N3929) );
  DFFPOSX1 \regZ_reg[6][4]  ( .D(n4901), .CLK(clk), .Q(N3925) );
  DFFPOSX1 \regZ_tri_enable_reg[6][4]  ( .D(n4900), .CLK(clk), .Q(N3926) );
  DFFPOSX1 \regZ_reg[6][5]  ( .D(n4899), .CLK(clk), .Q(N3922) );
  DFFPOSX1 \regZ_tri_enable_reg[6][5]  ( .D(n4898), .CLK(clk), .Q(N3923) );
  DFFPOSX1 \regZ_reg[6][6]  ( .D(n4897), .CLK(clk), .Q(N3919) );
  DFFPOSX1 \regZ_tri_enable_reg[6][6]  ( .D(n4896), .CLK(clk), .Q(N3920) );
  DFFPOSX1 \regZ_reg[6][7]  ( .D(n4895), .CLK(clk), .Q(N3916) );
  DFFPOSX1 \regZ_tri_enable_reg[6][7]  ( .D(n4894), .CLK(clk), .Q(N3917) );
  DFFPOSX1 \regZ_reg[7][0]  ( .D(n4893), .CLK(clk), .Q(N3961) );
  DFFPOSX1 \regZ_tri_enable_reg[7][0]  ( .D(n4892), .CLK(clk), .Q(N3962) );
  DFFPOSX1 \regZ_reg[7][1]  ( .D(n4891), .CLK(clk), .Q(N3958) );
  DFFPOSX1 \regZ_tri_enable_reg[7][1]  ( .D(n4890), .CLK(clk), .Q(N3959) );
  DFFPOSX1 \regZ_reg[7][2]  ( .D(n4889), .CLK(clk), .Q(N3955) );
  DFFPOSX1 \regZ_tri_enable_reg[7][2]  ( .D(n4888), .CLK(clk), .Q(N3956) );
  DFFPOSX1 \regZ_reg[7][3]  ( .D(n4887), .CLK(clk), .Q(N3952) );
  DFFPOSX1 \regZ_tri_enable_reg[7][3]  ( .D(n4886), .CLK(clk), .Q(N3953) );
  DFFPOSX1 \regZ_reg[7][4]  ( .D(n4885), .CLK(clk), .Q(N3949) );
  DFFPOSX1 \regZ_tri_enable_reg[7][4]  ( .D(n4884), .CLK(clk), .Q(N3950) );
  DFFPOSX1 \regZ_reg[7][5]  ( .D(n4883), .CLK(clk), .Q(N3946) );
  DFFPOSX1 \regZ_tri_enable_reg[7][5]  ( .D(n4882), .CLK(clk), .Q(N3947) );
  DFFPOSX1 \regZ_reg[7][6]  ( .D(n4881), .CLK(clk), .Q(N3943) );
  DFFPOSX1 \regZ_tri_enable_reg[7][6]  ( .D(n4880), .CLK(clk), .Q(N3944) );
  DFFPOSX1 \regZ_reg[7][7]  ( .D(n4879), .CLK(clk), .Q(N3940) );
  DFFPOSX1 \regZ_tri_enable_reg[7][7]  ( .D(n4878), .CLK(clk), .Q(N3941) );
  DFFPOSX1 \regZ_reg[8][0]  ( .D(n4877), .CLK(clk), .Q(N3985) );
  DFFPOSX1 \regZ_tri_enable_reg[8][0]  ( .D(n4876), .CLK(clk), .Q(N3986) );
  DFFPOSX1 \regZ_reg[8][1]  ( .D(n4875), .CLK(clk), .Q(N3982) );
  DFFPOSX1 \regZ_tri_enable_reg[8][1]  ( .D(n4874), .CLK(clk), .Q(N3983) );
  DFFPOSX1 \regZ_reg[8][2]  ( .D(n4873), .CLK(clk), .Q(N3979) );
  DFFPOSX1 \regZ_tri_enable_reg[8][2]  ( .D(n4872), .CLK(clk), .Q(N3980) );
  DFFPOSX1 \regZ_reg[8][3]  ( .D(n4871), .CLK(clk), .Q(N3976) );
  DFFPOSX1 \regZ_tri_enable_reg[8][3]  ( .D(n4870), .CLK(clk), .Q(N3977) );
  DFFPOSX1 \regZ_reg[8][4]  ( .D(n4869), .CLK(clk), .Q(N3973) );
  DFFPOSX1 \regZ_tri_enable_reg[8][4]  ( .D(n4868), .CLK(clk), .Q(N3974) );
  DFFPOSX1 \regZ_reg[8][5]  ( .D(n4867), .CLK(clk), .Q(N3970) );
  DFFPOSX1 \regZ_tri_enable_reg[8][5]  ( .D(n4866), .CLK(clk), .Q(N3971) );
  DFFPOSX1 \regZ_reg[8][6]  ( .D(n4865), .CLK(clk), .Q(N3967) );
  DFFPOSX1 \regZ_tri_enable_reg[8][6]  ( .D(n4864), .CLK(clk), .Q(N3968) );
  DFFPOSX1 \regZ_reg[8][7]  ( .D(n4863), .CLK(clk), .Q(N3964) );
  DFFPOSX1 \regZ_tri_enable_reg[8][7]  ( .D(n4862), .CLK(clk), .Q(N3965) );
  DFFPOSX1 \regZ_reg[9][0]  ( .D(n4861), .CLK(clk), .Q(N4009) );
  DFFPOSX1 \regZ_tri_enable_reg[9][0]  ( .D(n4860), .CLK(clk), .Q(N4010) );
  DFFPOSX1 \regZ_reg[9][1]  ( .D(n4859), .CLK(clk), .Q(N4006) );
  DFFPOSX1 \regZ_tri_enable_reg[9][1]  ( .D(n4858), .CLK(clk), .Q(N4007) );
  DFFPOSX1 \regZ_reg[9][2]  ( .D(n4857), .CLK(clk), .Q(N4003) );
  DFFPOSX1 \regZ_tri_enable_reg[9][2]  ( .D(n4856), .CLK(clk), .Q(N4004) );
  DFFPOSX1 \regZ_reg[9][3]  ( .D(n4855), .CLK(clk), .Q(N4000) );
  DFFPOSX1 \regZ_tri_enable_reg[9][3]  ( .D(n4854), .CLK(clk), .Q(N4001) );
  DFFPOSX1 \regZ_reg[9][4]  ( .D(n4853), .CLK(clk), .Q(N3997) );
  DFFPOSX1 \regZ_tri_enable_reg[9][4]  ( .D(n4852), .CLK(clk), .Q(N3998) );
  DFFPOSX1 \regZ_reg[9][5]  ( .D(n4851), .CLK(clk), .Q(N3994) );
  DFFPOSX1 \regZ_tri_enable_reg[9][5]  ( .D(n4850), .CLK(clk), .Q(N3995) );
  DFFPOSX1 \regZ_reg[9][6]  ( .D(n4849), .CLK(clk), .Q(N3991) );
  DFFPOSX1 \regZ_tri_enable_reg[9][6]  ( .D(n4848), .CLK(clk), .Q(N3992) );
  DFFPOSX1 \regZ_reg[9][7]  ( .D(n4847), .CLK(clk), .Q(N3988) );
  DFFPOSX1 \regZ_tri_enable_reg[9][7]  ( .D(n4846), .CLK(clk), .Q(N3989) );
  DFFPOSX1 \regZ_reg[16][0]  ( .D(n4845), .CLK(clk), .Q(N4177) );
  DFFPOSX1 \regZ_tri_enable_reg[16][0]  ( .D(n4844), .CLK(clk), .Q(N4178) );
  DFFPOSX1 \regZ_reg[16][1]  ( .D(n4843), .CLK(clk), .Q(N4174) );
  DFFPOSX1 \regZ_tri_enable_reg[16][1]  ( .D(n4842), .CLK(clk), .Q(N4175) );
  DFFPOSX1 \regZ_reg[16][2]  ( .D(n4841), .CLK(clk), .Q(N4171) );
  DFFPOSX1 \regZ_tri_enable_reg[16][2]  ( .D(n4840), .CLK(clk), .Q(N4172) );
  DFFPOSX1 \regZ_reg[16][3]  ( .D(n4839), .CLK(clk), .Q(N4168) );
  DFFPOSX1 \regZ_tri_enable_reg[16][3]  ( .D(n4838), .CLK(clk), .Q(N4169) );
  DFFPOSX1 \regZ_reg[16][4]  ( .D(n4837), .CLK(clk), .Q(N4165) );
  DFFPOSX1 \regZ_tri_enable_reg[16][4]  ( .D(n4836), .CLK(clk), .Q(N4166) );
  DFFPOSX1 \regZ_reg[16][5]  ( .D(n4835), .CLK(clk), .Q(N4162) );
  DFFPOSX1 \regZ_tri_enable_reg[16][5]  ( .D(n4834), .CLK(clk), .Q(N4163) );
  DFFPOSX1 \regZ_reg[16][6]  ( .D(n4833), .CLK(clk), .Q(N4159) );
  DFFPOSX1 \regZ_tri_enable_reg[16][6]  ( .D(n4832), .CLK(clk), .Q(N4160) );
  DFFPOSX1 \regZ_reg[16][7]  ( .D(n4831), .CLK(clk), .Q(N4156) );
  DFFPOSX1 \regZ_tri_enable_reg[16][7]  ( .D(n4830), .CLK(clk), .Q(N4157) );
  DFFPOSX1 \regZ_reg[17][0]  ( .D(n4829), .CLK(clk), .Q(N4201) );
  DFFPOSX1 \regZ_tri_enable_reg[17][0]  ( .D(n4828), .CLK(clk), .Q(N4202) );
  DFFPOSX1 \regZ_reg[17][1]  ( .D(n4827), .CLK(clk), .Q(N4198) );
  DFFPOSX1 \regZ_tri_enable_reg[17][1]  ( .D(n4826), .CLK(clk), .Q(N4199) );
  DFFPOSX1 \regZ_reg[17][2]  ( .D(n4825), .CLK(clk), .Q(N4195) );
  DFFPOSX1 \regZ_tri_enable_reg[17][2]  ( .D(n4824), .CLK(clk), .Q(N4196) );
  DFFPOSX1 \regZ_reg[17][3]  ( .D(n4823), .CLK(clk), .Q(N4192) );
  DFFPOSX1 \regZ_tri_enable_reg[17][3]  ( .D(n4822), .CLK(clk), .Q(N4193) );
  DFFPOSX1 \regZ_reg[17][4]  ( .D(n4821), .CLK(clk), .Q(N4189) );
  DFFPOSX1 \regZ_tri_enable_reg[17][4]  ( .D(n4820), .CLK(clk), .Q(N4190) );
  DFFPOSX1 \regZ_reg[17][5]  ( .D(n4819), .CLK(clk), .Q(N4186) );
  DFFPOSX1 \regZ_tri_enable_reg[17][5]  ( .D(n4818), .CLK(clk), .Q(N4187) );
  DFFPOSX1 \regZ_reg[17][6]  ( .D(n4817), .CLK(clk), .Q(N4183) );
  DFFPOSX1 \regZ_tri_enable_reg[17][6]  ( .D(n4816), .CLK(clk), .Q(N4184) );
  DFFPOSX1 \regZ_reg[17][7]  ( .D(n4815), .CLK(clk), .Q(N4180) );
  DFFPOSX1 \regZ_tri_enable_reg[17][7]  ( .D(n4814), .CLK(clk), .Q(N4181) );
  DFFPOSX1 \regZ_reg[24][0]  ( .D(n4813), .CLK(clk), .Q(N4369) );
  DFFPOSX1 \regZ_tri_enable_reg[24][0]  ( .D(n4812), .CLK(clk), .Q(N4370) );
  DFFPOSX1 \regZ_reg[24][1]  ( .D(n4811), .CLK(clk), .Q(N4366) );
  DFFPOSX1 \regZ_tri_enable_reg[24][1]  ( .D(n4810), .CLK(clk), .Q(N4367) );
  DFFPOSX1 \regZ_reg[24][2]  ( .D(n4809), .CLK(clk), .Q(N4363) );
  DFFPOSX1 \regZ_tri_enable_reg[24][2]  ( .D(n4808), .CLK(clk), .Q(N4364) );
  DFFPOSX1 \regZ_reg[24][3]  ( .D(n4807), .CLK(clk), .Q(N4360) );
  DFFPOSX1 \regZ_tri_enable_reg[24][3]  ( .D(n4806), .CLK(clk), .Q(N4361) );
  DFFPOSX1 \regZ_reg[24][4]  ( .D(n4805), .CLK(clk), .Q(N4357) );
  DFFPOSX1 \regZ_tri_enable_reg[24][4]  ( .D(n4804), .CLK(clk), .Q(N4358) );
  DFFPOSX1 \regZ_reg[24][5]  ( .D(n4803), .CLK(clk), .Q(N4354) );
  DFFPOSX1 \regZ_tri_enable_reg[24][5]  ( .D(n4802), .CLK(clk), .Q(N4355) );
  DFFPOSX1 \regZ_reg[24][6]  ( .D(n4801), .CLK(clk), .Q(N4351) );
  DFFPOSX1 \regZ_tri_enable_reg[24][6]  ( .D(n4800), .CLK(clk), .Q(N4352) );
  DFFPOSX1 \regZ_reg[24][7]  ( .D(n4799), .CLK(clk), .Q(N4348) );
  DFFPOSX1 \regZ_tri_enable_reg[24][7]  ( .D(n4798), .CLK(clk), .Q(N4349) );
  DFFPOSX1 \regZ_reg[14][0]  ( .D(n4797), .CLK(clk), .Q(N4129) );
  DFFPOSX1 \regZ_tri_enable_reg[14][0]  ( .D(n4796), .CLK(clk), .Q(N4130) );
  DFFPOSX1 \regZ_reg[14][1]  ( .D(n4795), .CLK(clk), .Q(N4126) );
  DFFPOSX1 \regZ_tri_enable_reg[14][1]  ( .D(n4794), .CLK(clk), .Q(N4127) );
  DFFPOSX1 \regZ_reg[14][2]  ( .D(n4793), .CLK(clk), .Q(N4123) );
  DFFPOSX1 \regZ_tri_enable_reg[14][2]  ( .D(n4792), .CLK(clk), .Q(N4124) );
  DFFPOSX1 \regZ_reg[14][3]  ( .D(n4791), .CLK(clk), .Q(N4120) );
  DFFPOSX1 \regZ_tri_enable_reg[14][3]  ( .D(n4790), .CLK(clk), .Q(N4121) );
  DFFPOSX1 \regZ_reg[14][4]  ( .D(n4789), .CLK(clk), .Q(N4117) );
  DFFPOSX1 \regZ_tri_enable_reg[14][4]  ( .D(n4788), .CLK(clk), .Q(N4118) );
  DFFPOSX1 \regZ_reg[14][5]  ( .D(n4787), .CLK(clk), .Q(N4114) );
  DFFPOSX1 \regZ_tri_enable_reg[14][5]  ( .D(n4786), .CLK(clk), .Q(N4115) );
  DFFPOSX1 \regZ_reg[14][6]  ( .D(n4785), .CLK(clk), .Q(N4111) );
  DFFPOSX1 \regZ_tri_enable_reg[14][6]  ( .D(n4784), .CLK(clk), .Q(N4112) );
  DFFPOSX1 \regZ_reg[14][7]  ( .D(n4783), .CLK(clk), .Q(N4108) );
  DFFPOSX1 \regZ_tri_enable_reg[14][7]  ( .D(n4782), .CLK(clk), .Q(N4109) );
  DFFPOSX1 \regZ_reg[15][0]  ( .D(n4781), .CLK(clk), .Q(N4153) );
  DFFPOSX1 \regZ_tri_enable_reg[15][0]  ( .D(n4780), .CLK(clk), .Q(N4154) );
  DFFPOSX1 \regZ_reg[15][1]  ( .D(n4779), .CLK(clk), .Q(N4150) );
  DFFPOSX1 \regZ_tri_enable_reg[15][1]  ( .D(n4778), .CLK(clk), .Q(N4151) );
  DFFPOSX1 \regZ_reg[15][2]  ( .D(n4777), .CLK(clk), .Q(N4147) );
  DFFPOSX1 \regZ_tri_enable_reg[15][2]  ( .D(n4776), .CLK(clk), .Q(N4148) );
  DFFPOSX1 \regZ_reg[15][3]  ( .D(n4775), .CLK(clk), .Q(N4144) );
  DFFPOSX1 \regZ_tri_enable_reg[15][3]  ( .D(n4774), .CLK(clk), .Q(N4145) );
  DFFPOSX1 \regZ_reg[15][4]  ( .D(n4773), .CLK(clk), .Q(N4141) );
  DFFPOSX1 \regZ_tri_enable_reg[15][4]  ( .D(n4772), .CLK(clk), .Q(N4142) );
  DFFPOSX1 \regZ_reg[15][5]  ( .D(n4771), .CLK(clk), .Q(N4138) );
  DFFPOSX1 \regZ_tri_enable_reg[15][5]  ( .D(n4770), .CLK(clk), .Q(N4139) );
  DFFPOSX1 \regZ_reg[15][6]  ( .D(n4769), .CLK(clk), .Q(N4135) );
  DFFPOSX1 \regZ_tri_enable_reg[15][6]  ( .D(n4768), .CLK(clk), .Q(N4136) );
  DFFPOSX1 \regZ_reg[15][7]  ( .D(n4767), .CLK(clk), .Q(N4132) );
  DFFPOSX1 \regZ_tri_enable_reg[15][7]  ( .D(n4766), .CLK(clk), .Q(N4133) );
  DFFPOSX1 \regZ_reg[22][0]  ( .D(n4765), .CLK(clk), .Q(N4321) );
  DFFPOSX1 \regZ_tri_enable_reg[22][0]  ( .D(n4764), .CLK(clk), .Q(N4322) );
  DFFPOSX1 \regZ_reg[22][1]  ( .D(n4763), .CLK(clk), .Q(N4318) );
  DFFPOSX1 \regZ_tri_enable_reg[22][1]  ( .D(n4762), .CLK(clk), .Q(N4319) );
  DFFPOSX1 \regZ_reg[22][2]  ( .D(n4761), .CLK(clk), .Q(N4315) );
  DFFPOSX1 \regZ_tri_enable_reg[22][2]  ( .D(n4760), .CLK(clk), .Q(N4316) );
  DFFPOSX1 \regZ_reg[22][3]  ( .D(n4759), .CLK(clk), .Q(N4312) );
  DFFPOSX1 \regZ_tri_enable_reg[22][3]  ( .D(n4758), .CLK(clk), .Q(N4313) );
  DFFPOSX1 \regZ_reg[22][4]  ( .D(n4757), .CLK(clk), .Q(N4309) );
  DFFPOSX1 \regZ_tri_enable_reg[22][4]  ( .D(n4756), .CLK(clk), .Q(N4310) );
  DFFPOSX1 \regZ_reg[22][5]  ( .D(n4755), .CLK(clk), .Q(N4306) );
  DFFPOSX1 \regZ_tri_enable_reg[22][5]  ( .D(n4754), .CLK(clk), .Q(N4307) );
  DFFPOSX1 \regZ_reg[22][6]  ( .D(n4753), .CLK(clk), .Q(N4303) );
  DFFPOSX1 \regZ_tri_enable_reg[22][6]  ( .D(n4752), .CLK(clk), .Q(N4304) );
  DFFPOSX1 \regZ_reg[22][7]  ( .D(n4751), .CLK(clk), .Q(N4300) );
  DFFPOSX1 \regZ_tri_enable_reg[22][7]  ( .D(n4750), .CLK(clk), .Q(N4301) );
  DFFPOSX1 \regZ_reg[23][0]  ( .D(n4749), .CLK(clk), .Q(N4345) );
  DFFPOSX1 \regZ_tri_enable_reg[23][0]  ( .D(n4748), .CLK(clk), .Q(N4346) );
  DFFPOSX1 \regZ_reg[23][1]  ( .D(n4747), .CLK(clk), .Q(N4342) );
  DFFPOSX1 \regZ_tri_enable_reg[23][1]  ( .D(n4746), .CLK(clk), .Q(N4343) );
  DFFPOSX1 \regZ_reg[23][2]  ( .D(n4745), .CLK(clk), .Q(N4339) );
  DFFPOSX1 \regZ_tri_enable_reg[23][2]  ( .D(n4744), .CLK(clk), .Q(N4340) );
  DFFPOSX1 \regZ_reg[23][3]  ( .D(n4743), .CLK(clk), .Q(N4336) );
  DFFPOSX1 \regZ_tri_enable_reg[23][3]  ( .D(n4742), .CLK(clk), .Q(N4337) );
  DFFPOSX1 \regZ_reg[23][4]  ( .D(n4741), .CLK(clk), .Q(N4333) );
  DFFPOSX1 \regZ_tri_enable_reg[23][4]  ( .D(n4740), .CLK(clk), .Q(N4334) );
  DFFPOSX1 \regZ_reg[23][5]  ( .D(n4739), .CLK(clk), .Q(N4330) );
  DFFPOSX1 \regZ_tri_enable_reg[23][5]  ( .D(n4738), .CLK(clk), .Q(N4331) );
  DFFPOSX1 \regZ_reg[23][6]  ( .D(n4737), .CLK(clk), .Q(N4327) );
  DFFPOSX1 \regZ_tri_enable_reg[23][6]  ( .D(n4736), .CLK(clk), .Q(N4328) );
  DFFPOSX1 \regZ_reg[23][7]  ( .D(n4735), .CLK(clk), .Q(N4324) );
  DFFPOSX1 \regZ_tri_enable_reg[23][7]  ( .D(n4734), .CLK(clk), .Q(N4325) );
  DFFPOSX1 \regZ_reg[13][0]  ( .D(n4733), .CLK(clk), .Q(N4105) );
  DFFPOSX1 \regZ_tri_enable_reg[13][0]  ( .D(n4732), .CLK(clk), .Q(N4106) );
  DFFPOSX1 \regZ_reg[13][1]  ( .D(n4731), .CLK(clk), .Q(N4102) );
  DFFPOSX1 \regZ_tri_enable_reg[13][1]  ( .D(n4730), .CLK(clk), .Q(N4103) );
  DFFPOSX1 \regZ_reg[13][2]  ( .D(n4729), .CLK(clk), .Q(N4099) );
  DFFPOSX1 \regZ_tri_enable_reg[13][2]  ( .D(n4728), .CLK(clk), .Q(N4100) );
  DFFPOSX1 \regZ_reg[13][3]  ( .D(n4727), .CLK(clk), .Q(N4096) );
  DFFPOSX1 \regZ_tri_enable_reg[13][3]  ( .D(n4726), .CLK(clk), .Q(N4097) );
  DFFPOSX1 \regZ_reg[13][4]  ( .D(n4725), .CLK(clk), .Q(N4093) );
  DFFPOSX1 \regZ_tri_enable_reg[13][4]  ( .D(n4724), .CLK(clk), .Q(N4094) );
  DFFPOSX1 \regZ_reg[13][5]  ( .D(n4723), .CLK(clk), .Q(N4090) );
  DFFPOSX1 \regZ_tri_enable_reg[13][5]  ( .D(n4722), .CLK(clk), .Q(N4091) );
  DFFPOSX1 \regZ_reg[13][6]  ( .D(n4721), .CLK(clk), .Q(N4087) );
  DFFPOSX1 \regZ_tri_enable_reg[13][6]  ( .D(n4720), .CLK(clk), .Q(N4088) );
  DFFPOSX1 \regZ_reg[13][7]  ( .D(n4719), .CLK(clk), .Q(N4084) );
  DFFPOSX1 \regZ_tri_enable_reg[13][7]  ( .D(n4718), .CLK(clk), .Q(N4085) );
  DFFPOSX1 \regZ_reg[20][0]  ( .D(n4717), .CLK(clk), .Q(N4273) );
  DFFPOSX1 \regZ_tri_enable_reg[20][0]  ( .D(n4716), .CLK(clk), .Q(N4274) );
  DFFPOSX1 \regZ_reg[20][1]  ( .D(n4715), .CLK(clk), .Q(N4270) );
  DFFPOSX1 \regZ_tri_enable_reg[20][1]  ( .D(n4714), .CLK(clk), .Q(N4271) );
  DFFPOSX1 \regZ_reg[20][2]  ( .D(n4713), .CLK(clk), .Q(N4267) );
  DFFPOSX1 \regZ_tri_enable_reg[20][2]  ( .D(n4712), .CLK(clk), .Q(N4268) );
  DFFPOSX1 \regZ_reg[20][3]  ( .D(n4711), .CLK(clk), .Q(N4264) );
  DFFPOSX1 \regZ_tri_enable_reg[20][3]  ( .D(n4710), .CLK(clk), .Q(N4265) );
  DFFPOSX1 \regZ_reg[20][4]  ( .D(n4709), .CLK(clk), .Q(N4261) );
  DFFPOSX1 \regZ_tri_enable_reg[20][4]  ( .D(n4708), .CLK(clk), .Q(N4262) );
  DFFPOSX1 \regZ_reg[20][5]  ( .D(n4707), .CLK(clk), .Q(N4258) );
  DFFPOSX1 \regZ_tri_enable_reg[20][5]  ( .D(n4706), .CLK(clk), .Q(N4259) );
  DFFPOSX1 \regZ_reg[20][6]  ( .D(n4705), .CLK(clk), .Q(N4255) );
  DFFPOSX1 \regZ_tri_enable_reg[20][6]  ( .D(n4704), .CLK(clk), .Q(N4256) );
  DFFPOSX1 \regZ_reg[20][7]  ( .D(n4703), .CLK(clk), .Q(N4252) );
  DFFPOSX1 \regZ_tri_enable_reg[20][7]  ( .D(n4702), .CLK(clk), .Q(N4253) );
  DFFPOSX1 \regZ_reg[21][0]  ( .D(n4701), .CLK(clk), .Q(N4297) );
  DFFPOSX1 \regZ_tri_enable_reg[21][0]  ( .D(n4700), .CLK(clk), .Q(N4298) );
  DFFPOSX1 \regZ_reg[21][1]  ( .D(n4699), .CLK(clk), .Q(N4294) );
  DFFPOSX1 \regZ_tri_enable_reg[21][1]  ( .D(n4698), .CLK(clk), .Q(N4295) );
  DFFPOSX1 \regZ_reg[21][2]  ( .D(n4697), .CLK(clk), .Q(N4291) );
  DFFPOSX1 \regZ_tri_enable_reg[21][2]  ( .D(n4696), .CLK(clk), .Q(N4292) );
  DFFPOSX1 \regZ_reg[21][3]  ( .D(n4695), .CLK(clk), .Q(N4288) );
  DFFPOSX1 \regZ_tri_enable_reg[21][3]  ( .D(n4694), .CLK(clk), .Q(N4289) );
  DFFPOSX1 \regZ_reg[21][4]  ( .D(n4693), .CLK(clk), .Q(N4285) );
  DFFPOSX1 \regZ_tri_enable_reg[21][4]  ( .D(n4692), .CLK(clk), .Q(N4286) );
  DFFPOSX1 \regZ_reg[21][5]  ( .D(n4691), .CLK(clk), .Q(N4282) );
  DFFPOSX1 \regZ_tri_enable_reg[21][5]  ( .D(n4690), .CLK(clk), .Q(N4283) );
  DFFPOSX1 \regZ_reg[21][6]  ( .D(n4689), .CLK(clk), .Q(N4279) );
  DFFPOSX1 \regZ_tri_enable_reg[21][6]  ( .D(n4688), .CLK(clk), .Q(N4280) );
  DFFPOSX1 \regZ_reg[21][7]  ( .D(n4687), .CLK(clk), .Q(N4276) );
  DFFPOSX1 \regZ_tri_enable_reg[21][7]  ( .D(n4686), .CLK(clk), .Q(N4277) );
  DFFPOSX1 \regZ_reg[10][0]  ( .D(n4685), .CLK(clk), .Q(N4033) );
  DFFPOSX1 \regZ_tri_enable_reg[10][0]  ( .D(n4684), .CLK(clk), .Q(N4034) );
  DFFPOSX1 \regZ_reg[10][1]  ( .D(n4683), .CLK(clk), .Q(N4030) );
  DFFPOSX1 \regZ_tri_enable_reg[10][1]  ( .D(n4682), .CLK(clk), .Q(N4031) );
  DFFPOSX1 \regZ_reg[10][2]  ( .D(n4681), .CLK(clk), .Q(N4027) );
  DFFPOSX1 \regZ_tri_enable_reg[10][2]  ( .D(n4680), .CLK(clk), .Q(N4028) );
  DFFPOSX1 \regZ_reg[10][3]  ( .D(n4679), .CLK(clk), .Q(N4024) );
  DFFPOSX1 \regZ_tri_enable_reg[10][3]  ( .D(n4678), .CLK(clk), .Q(N4025) );
  DFFPOSX1 \regZ_reg[10][4]  ( .D(n4677), .CLK(clk), .Q(N4021) );
  DFFPOSX1 \regZ_tri_enable_reg[10][4]  ( .D(n4676), .CLK(clk), .Q(N4022) );
  DFFPOSX1 \regZ_reg[10][5]  ( .D(n4675), .CLK(clk), .Q(N4018) );
  DFFPOSX1 \regZ_tri_enable_reg[10][5]  ( .D(n4674), .CLK(clk), .Q(N4019) );
  DFFPOSX1 \regZ_reg[10][6]  ( .D(n4673), .CLK(clk), .Q(N4015) );
  DFFPOSX1 \regZ_tri_enable_reg[10][6]  ( .D(n4672), .CLK(clk), .Q(N4016) );
  DFFPOSX1 \regZ_reg[10][7]  ( .D(n4671), .CLK(clk), .Q(N4012) );
  DFFPOSX1 \regZ_tri_enable_reg[10][7]  ( .D(n4670), .CLK(clk), .Q(N4013) );
  DFFPOSX1 \regZ_reg[11][0]  ( .D(n4669), .CLK(clk), .Q(N4057) );
  DFFPOSX1 \regZ_tri_enable_reg[11][0]  ( .D(n4668), .CLK(clk), .Q(N4058) );
  DFFPOSX1 \regZ_reg[11][1]  ( .D(n4667), .CLK(clk), .Q(N4054) );
  DFFPOSX1 \regZ_tri_enable_reg[11][1]  ( .D(n4666), .CLK(clk), .Q(N4055) );
  DFFPOSX1 \regZ_reg[11][2]  ( .D(n4665), .CLK(clk), .Q(N4051) );
  DFFPOSX1 \regZ_tri_enable_reg[11][2]  ( .D(n4664), .CLK(clk), .Q(N4052) );
  DFFPOSX1 \regZ_reg[11][3]  ( .D(n4663), .CLK(clk), .Q(N4048) );
  DFFPOSX1 \regZ_tri_enable_reg[11][3]  ( .D(n4662), .CLK(clk), .Q(N4049) );
  DFFPOSX1 \regZ_reg[11][4]  ( .D(n4661), .CLK(clk), .Q(N4045) );
  DFFPOSX1 \regZ_tri_enable_reg[11][4]  ( .D(n4660), .CLK(clk), .Q(N4046) );
  DFFPOSX1 \regZ_reg[11][5]  ( .D(n4659), .CLK(clk), .Q(N4042) );
  DFFPOSX1 \regZ_tri_enable_reg[11][5]  ( .D(n4658), .CLK(clk), .Q(N4043) );
  DFFPOSX1 \regZ_reg[11][6]  ( .D(n4657), .CLK(clk), .Q(N4039) );
  DFFPOSX1 \regZ_tri_enable_reg[11][6]  ( .D(n4656), .CLK(clk), .Q(N4040) );
  DFFPOSX1 \regZ_reg[11][7]  ( .D(n4655), .CLK(clk), .Q(N4036) );
  DFFPOSX1 \regZ_tri_enable_reg[11][7]  ( .D(n4654), .CLK(clk), .Q(N4037) );
  DFFPOSX1 \regZ_reg[18][0]  ( .D(n4653), .CLK(clk), .Q(N4225) );
  DFFPOSX1 \regZ_tri_enable_reg[18][0]  ( .D(n4652), .CLK(clk), .Q(N4226) );
  DFFPOSX1 \regZ_reg[18][1]  ( .D(n4651), .CLK(clk), .Q(N4222) );
  DFFPOSX1 \regZ_tri_enable_reg[18][1]  ( .D(n4650), .CLK(clk), .Q(N4223) );
  DFFPOSX1 \regZ_reg[18][2]  ( .D(n4649), .CLK(clk), .Q(N4219) );
  DFFPOSX1 \regZ_tri_enable_reg[18][2]  ( .D(n4648), .CLK(clk), .Q(N4220) );
  DFFPOSX1 \regZ_reg[18][3]  ( .D(n4647), .CLK(clk), .Q(N4216) );
  DFFPOSX1 \regZ_tri_enable_reg[18][3]  ( .D(n4646), .CLK(clk), .Q(N4217) );
  DFFPOSX1 \regZ_reg[18][4]  ( .D(n4645), .CLK(clk), .Q(N4213) );
  DFFPOSX1 \regZ_tri_enable_reg[18][4]  ( .D(n4644), .CLK(clk), .Q(N4214) );
  DFFPOSX1 \regZ_reg[18][5]  ( .D(n4643), .CLK(clk), .Q(N4210) );
  DFFPOSX1 \regZ_tri_enable_reg[18][5]  ( .D(n4642), .CLK(clk), .Q(N4211) );
  DFFPOSX1 \regZ_reg[18][6]  ( .D(n4641), .CLK(clk), .Q(N4207) );
  DFFPOSX1 \regZ_tri_enable_reg[18][6]  ( .D(n4640), .CLK(clk), .Q(N4208) );
  DFFPOSX1 \regZ_reg[18][7]  ( .D(n4639), .CLK(clk), .Q(N4204) );
  DFFPOSX1 \regZ_tri_enable_reg[18][7]  ( .D(n4638), .CLK(clk), .Q(N4205) );
  DFFPOSX1 \regZ_reg[19][0]  ( .D(n4637), .CLK(clk), .Q(N4249) );
  DFFPOSX1 \regZ_tri_enable_reg[19][0]  ( .D(n4636), .CLK(clk), .Q(N4250) );
  DFFPOSX1 \regZ_reg[19][1]  ( .D(n4635), .CLK(clk), .Q(N4246) );
  DFFPOSX1 \regZ_tri_enable_reg[19][1]  ( .D(n4634), .CLK(clk), .Q(N4247) );
  DFFPOSX1 \regZ_reg[19][2]  ( .D(n4633), .CLK(clk), .Q(N4243) );
  DFFPOSX1 \regZ_tri_enable_reg[19][2]  ( .D(n4632), .CLK(clk), .Q(N4244) );
  DFFPOSX1 \regZ_reg[19][3]  ( .D(n4631), .CLK(clk), .Q(N4240) );
  DFFPOSX1 \regZ_tri_enable_reg[19][3]  ( .D(n4630), .CLK(clk), .Q(N4241) );
  DFFPOSX1 \regZ_reg[19][4]  ( .D(n4629), .CLK(clk), .Q(N4237) );
  DFFPOSX1 \regZ_tri_enable_reg[19][4]  ( .D(n4628), .CLK(clk), .Q(N4238) );
  DFFPOSX1 \regZ_reg[19][5]  ( .D(n4627), .CLK(clk), .Q(N4234) );
  DFFPOSX1 \regZ_tri_enable_reg[19][5]  ( .D(n4626), .CLK(clk), .Q(N4235) );
  DFFPOSX1 \regZ_reg[19][6]  ( .D(n4625), .CLK(clk), .Q(N4231) );
  DFFPOSX1 \regZ_tri_enable_reg[19][6]  ( .D(n4624), .CLK(clk), .Q(N4232) );
  DFFPOSX1 \regZ_reg[19][7]  ( .D(n4623), .CLK(clk), .Q(N4228) );
  DFFPOSX1 \regZ_tri_enable_reg[19][7]  ( .D(n4622), .CLK(clk), .Q(N4229) );
  DFFPOSX1 \regZ_tri_enable_reg[2][7]  ( .D(n4621), .CLK(clk), .Q(N3821) );
  DFFPOSX1 \regZ_reg[2][7]  ( .D(n4620), .CLK(clk), .Q(N3820) );
  DFFPOSX1 \regZ_tri_enable_reg[2][6]  ( .D(n4619), .CLK(clk), .Q(N3824) );
  DFFPOSX1 \regZ_reg[2][6]  ( .D(n4618), .CLK(clk), .Q(N3823) );
  DFFPOSX1 \regZ_tri_enable_reg[2][5]  ( .D(n4617), .CLK(clk), .Q(N3827) );
  DFFPOSX1 \regZ_reg[2][5]  ( .D(n4616), .CLK(clk), .Q(N3826) );
  DFFPOSX1 \regZ_tri_enable_reg[2][4]  ( .D(n4615), .CLK(clk), .Q(N3830) );
  DFFPOSX1 \regZ_reg[2][4]  ( .D(n4614), .CLK(clk), .Q(N3829) );
  DFFPOSX1 \regZ_tri_enable_reg[2][3]  ( .D(n4613), .CLK(clk), .Q(N3833) );
  DFFPOSX1 \regZ_reg[2][3]  ( .D(n4612), .CLK(clk), .Q(N3832) );
  DFFPOSX1 \regZ_tri_enable_reg[2][2]  ( .D(n4611), .CLK(clk), .Q(N3836) );
  DFFPOSX1 \regZ_reg[2][2]  ( .D(n4610), .CLK(clk), .Q(N3835) );
  DFFPOSX1 \regZ_tri_enable_reg[2][1]  ( .D(n4609), .CLK(clk), .Q(N3839) );
  DFFPOSX1 \regZ_reg[2][1]  ( .D(n4608), .CLK(clk), .Q(N3838) );
  DFFPOSX1 \regZ_tri_enable_reg[2][0]  ( .D(n4607), .CLK(clk), .Q(N3842) );
  DFFPOSX1 \regZ_reg[2][0]  ( .D(n4606), .CLK(clk), .Q(N3841) );
  DFFPOSX1 \regZ_tri_enable_reg[1][7]  ( .D(n4605), .CLK(clk), .Q(N3797) );
  DFFPOSX1 \regZ_reg[1][7]  ( .D(n4604), .CLK(clk), .Q(N3796) );
  DFFPOSX1 \regZ_tri_enable_reg[1][6]  ( .D(n4603), .CLK(clk), .Q(N3800) );
  DFFPOSX1 \regZ_reg[1][6]  ( .D(n4602), .CLK(clk), .Q(N3799) );
  DFFPOSX1 \regZ_tri_enable_reg[1][5]  ( .D(n4601), .CLK(clk), .Q(N3803) );
  DFFPOSX1 \regZ_reg[1][5]  ( .D(n4600), .CLK(clk), .Q(N3802) );
  DFFPOSX1 \regZ_tri_enable_reg[1][4]  ( .D(n4599), .CLK(clk), .Q(N3806) );
  DFFPOSX1 \regZ_reg[1][4]  ( .D(n4598), .CLK(clk), .Q(N3805) );
  DFFPOSX1 \regZ_tri_enable_reg[1][3]  ( .D(n4597), .CLK(clk), .Q(N3809) );
  DFFPOSX1 \regZ_reg[1][3]  ( .D(n4596), .CLK(clk), .Q(N3808) );
  DFFPOSX1 \regZ_tri_enable_reg[1][2]  ( .D(n4595), .CLK(clk), .Q(N3812) );
  DFFPOSX1 \regZ_reg[1][2]  ( .D(n4594), .CLK(clk), .Q(N3811) );
  DFFPOSX1 \regZ_tri_enable_reg[1][1]  ( .D(n4593), .CLK(clk), .Q(N3815) );
  DFFPOSX1 \regZ_reg[1][1]  ( .D(n4592), .CLK(clk), .Q(N3814) );
  DFFPOSX1 \regZ_tri_enable_reg[1][0]  ( .D(n4591), .CLK(clk), .Q(N3818) );
  DFFPOSX1 \regZ_reg[1][0]  ( .D(n4590), .CLK(clk), .Q(N3817) );
  DFFPOSX1 \Out_bThres_reg[0]  ( .D(n4589), .CLK(clk), .Q(\Out_bThres[0] ) );
  DFFPOSX1 \tpSum_reg[7]  ( .D(n4588), .CLK(clk), .Q(tpSum[7]) );
  DFFPOSX1 \tpSum_reg[8]  ( .D(n4587), .CLK(clk), .Q(tpSum[8]) );
  DFFPOSX1 \tpSum_reg[9]  ( .D(n4586), .CLK(clk), .Q(tpSum[9]) );
  DFFPOSX1 \tpSum_reg[10]  ( .D(n4585), .CLK(clk), .Q(tpSum[10]) );
  DFFPOSX1 \tpSum_reg[11]  ( .D(n4584), .CLK(clk), .Q(tpSum[11]) );
  DFFPOSX1 \tpSum_reg[12]  ( .D(n4583), .CLK(clk), .Q(tpSum[12]) );
  DFFPOSX1 \tpSum_reg[13]  ( .D(n4582), .CLK(clk), .Q(tpSum[13]) );
  DFFPOSX1 \tpSum_reg[14]  ( .D(n4581), .CLK(clk), .Q(tpSum[14]) );
  DFFPOSX1 \Out_gf_reg[7]  ( .D(n8315), .CLK(clk), .Q(Out_gf[7]) );
  DFFPOSX1 \OutData_reg[7]  ( .D(n4579), .CLK(clk), .Q(N4468) );
  DFFPOSX1 \Out_gf_reg[6]  ( .D(n8316), .CLK(clk), .Q(Out_gf[6]) );
  DFFPOSX1 \OutData_reg[6]  ( .D(n4577), .CLK(clk), .Q(N4471) );
  DFFPOSX1 \Out_gf_reg[5]  ( .D(n8317), .CLK(clk), .Q(Out_gf[5]) );
  DFFPOSX1 \OutData_reg[5]  ( .D(n4575), .CLK(clk), .Q(N4474) );
  DFFPOSX1 \Out_gf_reg[4]  ( .D(n8318), .CLK(clk), .Q(Out_gf[4]) );
  DFFPOSX1 \OutData_reg[4]  ( .D(n4573), .CLK(clk), .Q(N4477) );
  DFFPOSX1 \Out_gf_reg[3]  ( .D(n8319), .CLK(clk), .Q(Out_gf[3]) );
  DFFPOSX1 \OutData_reg[3]  ( .D(n4571), .CLK(clk), .Q(N4480) );
  DFFPOSX1 \Out_gf_reg[2]  ( .D(n8320), .CLK(clk), .Q(Out_gf[2]) );
  DFFPOSX1 \OutData_reg[2]  ( .D(n4569), .CLK(clk), .Q(N4483) );
  DFFPOSX1 \Out_gf_reg[1]  ( .D(n8321), .CLK(clk), .Q(Out_gf[1]) );
  DFFPOSX1 \OutData_reg[1]  ( .D(n4567), .CLK(clk), .Q(N4486) );
  DFFPOSX1 \Out_gf_reg[0]  ( .D(n8322), .CLK(clk), .Q(Out_gf[0]) );
  DFFPOSX1 \OutData_reg[0]  ( .D(n4565), .CLK(clk), .Q(N4489) );
  TBUFX1 \dx_tri[0]  ( .A(n15427), .EN(n15394), .Y(dx[0]) );
  TBUFX1 \dy_tri[0]  ( .A(n15428), .EN(n15429), .Y(dy[0]) );
  TBUFX1 \OutData_tri[0]  ( .A(n15853), .EN(n15322), .Y(OutData[0]) );
  TBUFX1 \OutData_tri[1]  ( .A(n15852), .EN(n15321), .Y(OutData[1]) );
  TBUFX1 \OutData_tri[2]  ( .A(n15851), .EN(n15320), .Y(OutData[2]) );
  TBUFX1 \OutData_tri[3]  ( .A(n15850), .EN(n15319), .Y(OutData[3]) );
  TBUFX1 \OutData_tri[4]  ( .A(n15849), .EN(n15318), .Y(OutData[4]) );
  TBUFX1 \OutData_tri[5]  ( .A(n15848), .EN(n15317), .Y(OutData[5]) );
  TBUFX1 \OutData_tri[6]  ( .A(n15847), .EN(n15316), .Y(OutData[6]) );
  TBUFX1 \OutData_tri[7]  ( .A(n15846), .EN(n15315), .Y(OutData[7]) );
  TBUFX1 \fGy_tri[0]  ( .A(n15438), .EN(n15378), .Y(fGy[0]) );
  TBUFX1 \fGy_tri[1]  ( .A(n15439), .EN(n15379), .Y(fGy[1]) );
  TBUFX1 \fGy_tri[2]  ( .A(n15440), .EN(n15380), .Y(fGy[2]) );
  TBUFX1 \fGy_tri[3]  ( .A(n15441), .EN(n15381), .Y(fGy[3]) );
  TBUFX1 \fGy_tri[4]  ( .A(n15442), .EN(n15382), .Y(fGy[4]) );
  TBUFX1 \fGy_tri[5]  ( .A(n15443), .EN(n15383), .Y(fGy[5]) );
  TBUFX1 \fGy_tri[6]  ( .A(n15444), .EN(n15384), .Y(fGy[6]) );
  TBUFX1 \fGy_tri[7]  ( .A(n15445), .EN(n15385), .Y(fGy[7]) );
  TBUFX1 \Out_direction_tri[0]  ( .A(n15462), .EN(n15463), .Y(Out_direction[0]) );
  TBUFX1 \Out_direction_tri[1]  ( .A(n15464), .EN(n15465), .Y(Out_direction[1]) );
  TBUFX1 \Out_direction_tri[2]  ( .A(n15466), .EN(n15467), .Y(Out_direction[2]) );
  TBUFX1 \Out_direction_tri[3]  ( .A(n15468), .EN(n15469), .Y(Out_direction[3]) );
  TBUFX1 \Out_direction_tri[4]  ( .A(n15470), .EN(n15471), .Y(Out_direction[4]) );
  TBUFX1 \Out_direction_tri[5]  ( .A(n15472), .EN(n15473), .Y(Out_direction[5]) );
  TBUFX1 \Out_direction_tri[6]  ( .A(n15474), .EN(n15475), .Y(Out_direction[6]) );
  TBUFX1 \Out_direction_tri[7]  ( .A(n15476), .EN(n15477), .Y(Out_direction[7]) );
  TBUFX1 \Out_gradient_tri[0]  ( .A(n15454), .EN(n15430), .Y(Out_gradient[0])
         );
  TBUFX1 \Out_gradient_tri[1]  ( .A(n15455), .EN(n15431), .Y(Out_gradient[1])
         );
  TBUFX1 \Out_gradient_tri[2]  ( .A(n15456), .EN(n15432), .Y(Out_gradient[2])
         );
  TBUFX1 \Out_gradient_tri[3]  ( .A(n15457), .EN(n15433), .Y(Out_gradient[3])
         );
  TBUFX1 \Out_gradient_tri[4]  ( .A(n15458), .EN(n15434), .Y(Out_gradient[4])
         );
  TBUFX1 \Out_gradient_tri[5]  ( .A(n15459), .EN(n15435), .Y(Out_gradient[5])
         );
  TBUFX1 \Out_gradient_tri[6]  ( .A(n15460), .EN(n15436), .Y(Out_gradient[6])
         );
  TBUFX1 \Out_gradient_tri[7]  ( .A(n15461), .EN(n15437), .Y(Out_gradient[7])
         );
  TBUFX1 \fGx_tri[0]  ( .A(n15446), .EN(n15393), .Y(fGx[0]) );
  TBUFX1 \fGx_tri[1]  ( .A(n15447), .EN(n15392), .Y(fGx[1]) );
  TBUFX1 \fGx_tri[2]  ( .A(n15448), .EN(n15391), .Y(fGx[2]) );
  TBUFX1 \fGx_tri[3]  ( .A(n15449), .EN(n15390), .Y(fGx[3]) );
  TBUFX1 \fGx_tri[4]  ( .A(n15450), .EN(n15389), .Y(fGx[4]) );
  TBUFX1 \fGx_tri[5]  ( .A(n15451), .EN(n15388), .Y(fGx[5]) );
  TBUFX1 \fGx_tri[6]  ( .A(n15452), .EN(n15387), .Y(fGx[6]) );
  TBUFX1 \fGx_tri[7]  ( .A(n15453), .EN(n15386), .Y(fGx[7]) );
  TBUFX1 \regZ_tri[24][0]  ( .A(n15622), .EN(n15623), .Y(\regZ[24][0] ) );
  TBUFX1 \regZ_tri[24][1]  ( .A(n15624), .EN(n15625), .Y(\regZ[24][1] ) );
  TBUFX1 \regZ_tri[24][2]  ( .A(n15626), .EN(n15627), .Y(\regZ[24][2] ) );
  TBUFX1 \regZ_tri[24][3]  ( .A(n15628), .EN(n15629), .Y(\regZ[24][3] ) );
  TBUFX1 \regZ_tri[24][4]  ( .A(n15630), .EN(n15631), .Y(\regZ[24][4] ) );
  TBUFX1 \regZ_tri[24][5]  ( .A(n15632), .EN(n15633), .Y(\regZ[24][5] ) );
  TBUFX1 \regZ_tri[24][6]  ( .A(n15634), .EN(n15635), .Y(\regZ[24][6] ) );
  TBUFX1 \regZ_tri[24][7]  ( .A(n15636), .EN(n15637), .Y(\regZ[24][7] ) );
  TBUFX1 \regZ_tri[23][0]  ( .A(n15686), .EN(n15687), .Y(\regZ[23][0] ) );
  TBUFX1 \regZ_tri[23][1]  ( .A(n15688), .EN(n15689), .Y(\regZ[23][1] ) );
  TBUFX1 \regZ_tri[23][2]  ( .A(n15690), .EN(n15691), .Y(\regZ[23][2] ) );
  TBUFX1 \regZ_tri[23][3]  ( .A(n15692), .EN(n15693), .Y(\regZ[23][3] ) );
  TBUFX1 \regZ_tri[23][4]  ( .A(n15694), .EN(n15695), .Y(\regZ[23][4] ) );
  TBUFX1 \regZ_tri[23][5]  ( .A(n15696), .EN(n15697), .Y(\regZ[23][5] ) );
  TBUFX1 \regZ_tri[23][6]  ( .A(n15698), .EN(n15699), .Y(\regZ[23][6] ) );
  TBUFX1 \regZ_tri[23][7]  ( .A(n15700), .EN(n15701), .Y(\regZ[23][7] ) );
  TBUFX1 \regZ_tri[22][0]  ( .A(n15670), .EN(n15671), .Y(\regZ[22][0] ) );
  TBUFX1 \regZ_tri[22][1]  ( .A(n15672), .EN(n15673), .Y(\regZ[22][1] ) );
  TBUFX1 \regZ_tri[22][2]  ( .A(n15674), .EN(n15675), .Y(\regZ[22][2] ) );
  TBUFX1 \regZ_tri[22][3]  ( .A(n15676), .EN(n15677), .Y(\regZ[22][3] ) );
  TBUFX1 \regZ_tri[22][4]  ( .A(n15678), .EN(n15679), .Y(\regZ[22][4] ) );
  TBUFX1 \regZ_tri[22][5]  ( .A(n15680), .EN(n15681), .Y(\regZ[22][5] ) );
  TBUFX1 \regZ_tri[22][6]  ( .A(n15682), .EN(n15683), .Y(\regZ[22][6] ) );
  TBUFX1 \regZ_tri[22][7]  ( .A(n15684), .EN(n15685), .Y(\regZ[22][7] ) );
  TBUFX1 \regZ_tri[21][0]  ( .A(n15734), .EN(n15735), .Y(\regZ[21][0] ) );
  TBUFX1 \regZ_tri[21][1]  ( .A(n15736), .EN(n15737), .Y(\regZ[21][1] ) );
  TBUFX1 \regZ_tri[21][2]  ( .A(n15738), .EN(n15739), .Y(\regZ[21][2] ) );
  TBUFX1 \regZ_tri[21][3]  ( .A(n15740), .EN(n15741), .Y(\regZ[21][3] ) );
  TBUFX1 \regZ_tri[21][4]  ( .A(n15742), .EN(n15743), .Y(\regZ[21][4] ) );
  TBUFX1 \regZ_tri[21][5]  ( .A(n15744), .EN(n15745), .Y(\regZ[21][5] ) );
  TBUFX1 \regZ_tri[21][6]  ( .A(n15746), .EN(n15747), .Y(\regZ[21][6] ) );
  TBUFX1 \regZ_tri[21][7]  ( .A(n15748), .EN(n15749), .Y(\regZ[21][7] ) );
  TBUFX1 \regZ_tri[20][0]  ( .A(n15718), .EN(n15719), .Y(\regZ[20][0] ) );
  TBUFX1 \regZ_tri[20][1]  ( .A(n15720), .EN(n15721), .Y(\regZ[20][1] ) );
  TBUFX1 \regZ_tri[20][2]  ( .A(n15722), .EN(n15723), .Y(\regZ[20][2] ) );
  TBUFX1 \regZ_tri[20][3]  ( .A(n15724), .EN(n15725), .Y(\regZ[20][3] ) );
  TBUFX1 \regZ_tri[20][4]  ( .A(n15726), .EN(n15727), .Y(\regZ[20][4] ) );
  TBUFX1 \regZ_tri[20][5]  ( .A(n15728), .EN(n15729), .Y(\regZ[20][5] ) );
  TBUFX1 \regZ_tri[20][6]  ( .A(n15730), .EN(n15731), .Y(\regZ[20][6] ) );
  TBUFX1 \regZ_tri[20][7]  ( .A(n15732), .EN(n15733), .Y(\regZ[20][7] ) );
  TBUFX1 \regZ_tri[19][0]  ( .A(n15798), .EN(n15799), .Y(\regZ[19][0] ) );
  TBUFX1 \regZ_tri[19][1]  ( .A(n15800), .EN(n15801), .Y(\regZ[19][1] ) );
  TBUFX1 \regZ_tri[19][2]  ( .A(n15802), .EN(n15803), .Y(\regZ[19][2] ) );
  TBUFX1 \regZ_tri[19][3]  ( .A(n15804), .EN(n15805), .Y(\regZ[19][3] ) );
  TBUFX1 \regZ_tri[19][4]  ( .A(n15806), .EN(n15807), .Y(\regZ[19][4] ) );
  TBUFX1 \regZ_tri[19][5]  ( .A(n15808), .EN(n15809), .Y(\regZ[19][5] ) );
  TBUFX1 \regZ_tri[19][6]  ( .A(n15810), .EN(n15811), .Y(\regZ[19][6] ) );
  TBUFX1 \regZ_tri[19][7]  ( .A(n15812), .EN(n15813), .Y(\regZ[19][7] ) );
  TBUFX1 \regZ_tri[18][0]  ( .A(n15782), .EN(n15783), .Y(\regZ[18][0] ) );
  TBUFX1 \regZ_tri[18][1]  ( .A(n15784), .EN(n15785), .Y(\regZ[18][1] ) );
  TBUFX1 \regZ_tri[18][2]  ( .A(n15786), .EN(n15787), .Y(\regZ[18][2] ) );
  TBUFX1 \regZ_tri[18][3]  ( .A(n15788), .EN(n15789), .Y(\regZ[18][3] ) );
  TBUFX1 \regZ_tri[18][4]  ( .A(n15790), .EN(n15791), .Y(\regZ[18][4] ) );
  TBUFX1 \regZ_tri[18][5]  ( .A(n15792), .EN(n15793), .Y(\regZ[18][5] ) );
  TBUFX1 \regZ_tri[18][6]  ( .A(n15794), .EN(n15795), .Y(\regZ[18][6] ) );
  TBUFX1 \regZ_tri[18][7]  ( .A(n15796), .EN(n15797), .Y(\regZ[18][7] ) );
  TBUFX1 \regZ_tri[17][0]  ( .A(n15606), .EN(n15607), .Y(\regZ[17][0] ) );
  TBUFX1 \regZ_tri[17][1]  ( .A(n15608), .EN(n15609), .Y(\regZ[17][1] ) );
  TBUFX1 \regZ_tri[17][2]  ( .A(n15610), .EN(n15611), .Y(\regZ[17][2] ) );
  TBUFX1 \regZ_tri[17][3]  ( .A(n15612), .EN(n15613), .Y(\regZ[17][3] ) );
  TBUFX1 \regZ_tri[17][4]  ( .A(n15614), .EN(n15615), .Y(\regZ[17][4] ) );
  TBUFX1 \regZ_tri[17][5]  ( .A(n15616), .EN(n15617), .Y(\regZ[17][5] ) );
  TBUFX1 \regZ_tri[17][6]  ( .A(n15618), .EN(n15619), .Y(\regZ[17][6] ) );
  TBUFX1 \regZ_tri[17][7]  ( .A(n15620), .EN(n15621), .Y(\regZ[17][7] ) );
  TBUFX1 \regZ_tri[16][0]  ( .A(n15590), .EN(n15591), .Y(\regZ[16][0] ) );
  TBUFX1 \regZ_tri[16][1]  ( .A(n15592), .EN(n15593), .Y(\regZ[16][1] ) );
  TBUFX1 \regZ_tri[16][2]  ( .A(n15594), .EN(n15595), .Y(\regZ[16][2] ) );
  TBUFX1 \regZ_tri[16][3]  ( .A(n15596), .EN(n15597), .Y(\regZ[16][3] ) );
  TBUFX1 \regZ_tri[16][4]  ( .A(n15598), .EN(n15599), .Y(\regZ[16][4] ) );
  TBUFX1 \regZ_tri[16][5]  ( .A(n15600), .EN(n15601), .Y(\regZ[16][5] ) );
  TBUFX1 \regZ_tri[16][6]  ( .A(n15602), .EN(n15603), .Y(\regZ[16][6] ) );
  TBUFX1 \regZ_tri[16][7]  ( .A(n15604), .EN(n15605), .Y(\regZ[16][7] ) );
  TBUFX1 \regZ_tri[15][0]  ( .A(n15654), .EN(n15655), .Y(\regZ[15][0] ) );
  TBUFX1 \regZ_tri[15][1]  ( .A(n15656), .EN(n15657), .Y(\regZ[15][1] ) );
  TBUFX1 \regZ_tri[15][2]  ( .A(n15658), .EN(n15659), .Y(\regZ[15][2] ) );
  TBUFX1 \regZ_tri[15][3]  ( .A(n15660), .EN(n15661), .Y(\regZ[15][3] ) );
  TBUFX1 \regZ_tri[15][4]  ( .A(n15662), .EN(n15663), .Y(\regZ[15][4] ) );
  TBUFX1 \regZ_tri[15][5]  ( .A(n15664), .EN(n15665), .Y(\regZ[15][5] ) );
  TBUFX1 \regZ_tri[15][6]  ( .A(n15666), .EN(n15667), .Y(\regZ[15][6] ) );
  TBUFX1 \regZ_tri[15][7]  ( .A(n15668), .EN(n15669), .Y(\regZ[15][7] ) );
  TBUFX1 \regZ_tri[14][0]  ( .A(n15638), .EN(n15639), .Y(\regZ[14][0] ) );
  TBUFX1 \regZ_tri[14][1]  ( .A(n15640), .EN(n15641), .Y(\regZ[14][1] ) );
  TBUFX1 \regZ_tri[14][2]  ( .A(n15642), .EN(n15643), .Y(\regZ[14][2] ) );
  TBUFX1 \regZ_tri[14][3]  ( .A(n15644), .EN(n15645), .Y(\regZ[14][3] ) );
  TBUFX1 \regZ_tri[14][4]  ( .A(n15646), .EN(n15647), .Y(\regZ[14][4] ) );
  TBUFX1 \regZ_tri[14][5]  ( .A(n15648), .EN(n15649), .Y(\regZ[14][5] ) );
  TBUFX1 \regZ_tri[14][6]  ( .A(n15650), .EN(n15651), .Y(\regZ[14][6] ) );
  TBUFX1 \regZ_tri[14][7]  ( .A(n15652), .EN(n15653), .Y(\regZ[14][7] ) );
  TBUFX1 \regZ_tri[13][0]  ( .A(n15702), .EN(n15703), .Y(\regZ[13][0] ) );
  TBUFX1 \regZ_tri[13][1]  ( .A(n15704), .EN(n15705), .Y(\regZ[13][1] ) );
  TBUFX1 \regZ_tri[13][2]  ( .A(n15706), .EN(n15707), .Y(\regZ[13][2] ) );
  TBUFX1 \regZ_tri[13][3]  ( .A(n15708), .EN(n15709), .Y(\regZ[13][3] ) );
  TBUFX1 \regZ_tri[13][4]  ( .A(n15710), .EN(n15711), .Y(\regZ[13][4] ) );
  TBUFX1 \regZ_tri[13][5]  ( .A(n15712), .EN(n15713), .Y(\regZ[13][5] ) );
  TBUFX1 \regZ_tri[13][6]  ( .A(n15714), .EN(n15715), .Y(\regZ[13][6] ) );
  TBUFX1 \regZ_tri[13][7]  ( .A(n15716), .EN(n15717), .Y(\regZ[13][7] ) );
  TBUFX1 \regZ_tri[12][0]  ( .A(n15395), .EN(n15396), .Y(\regZ[12][0] ) );
  TBUFX1 \regZ_tri[12][1]  ( .A(n15410), .EN(n15409), .Y(\regZ[12][1] ) );
  TBUFX1 \regZ_tri[12][2]  ( .A(n15408), .EN(n15407), .Y(\regZ[12][2] ) );
  TBUFX1 \regZ_tri[12][3]  ( .A(n15406), .EN(n15405), .Y(\regZ[12][3] ) );
  TBUFX1 \regZ_tri[12][4]  ( .A(n15404), .EN(n15403), .Y(\regZ[12][4] ) );
  TBUFX1 \regZ_tri[12][5]  ( .A(n15402), .EN(n15401), .Y(\regZ[12][5] ) );
  TBUFX1 \regZ_tri[12][6]  ( .A(n15400), .EN(n15399), .Y(\regZ[12][6] ) );
  TBUFX1 \regZ_tri[12][7]  ( .A(n15398), .EN(n15397), .Y(\regZ[12][7] ) );
  TBUFX1 \regZ_tri[11][0]  ( .A(n15766), .EN(n15767), .Y(\regZ[11][0] ) );
  TBUFX1 \regZ_tri[11][1]  ( .A(n15768), .EN(n15769), .Y(\regZ[11][1] ) );
  TBUFX1 \regZ_tri[11][2]  ( .A(n15770), .EN(n15771), .Y(\regZ[11][2] ) );
  TBUFX1 \regZ_tri[11][3]  ( .A(n15772), .EN(n15773), .Y(\regZ[11][3] ) );
  TBUFX1 \regZ_tri[11][4]  ( .A(n15774), .EN(n15775), .Y(\regZ[11][4] ) );
  TBUFX1 \regZ_tri[11][5]  ( .A(n15776), .EN(n15777), .Y(\regZ[11][5] ) );
  TBUFX1 \regZ_tri[11][6]  ( .A(n15778), .EN(n15779), .Y(\regZ[11][6] ) );
  TBUFX1 \regZ_tri[11][7]  ( .A(n15780), .EN(n15781), .Y(\regZ[11][7] ) );
  TBUFX1 \regZ_tri[10][0]  ( .A(n15750), .EN(n15751), .Y(\regZ[10][0] ) );
  TBUFX1 \regZ_tri[10][1]  ( .A(n15752), .EN(n15753), .Y(\regZ[10][1] ) );
  TBUFX1 \regZ_tri[10][2]  ( .A(n15754), .EN(n15755), .Y(\regZ[10][2] ) );
  TBUFX1 \regZ_tri[10][3]  ( .A(n15756), .EN(n15757), .Y(\regZ[10][3] ) );
  TBUFX1 \regZ_tri[10][4]  ( .A(n15758), .EN(n15759), .Y(\regZ[10][4] ) );
  TBUFX1 \regZ_tri[10][5]  ( .A(n15760), .EN(n15761), .Y(\regZ[10][5] ) );
  TBUFX1 \regZ_tri[10][6]  ( .A(n15762), .EN(n15763), .Y(\regZ[10][6] ) );
  TBUFX1 \regZ_tri[10][7]  ( .A(n15764), .EN(n15765), .Y(\regZ[10][7] ) );
  TBUFX1 \regZ_tri[9][0]  ( .A(n15574), .EN(n15575), .Y(\regZ[9][0] ) );
  TBUFX1 \regZ_tri[9][1]  ( .A(n15576), .EN(n15577), .Y(\regZ[9][1] ) );
  TBUFX1 \regZ_tri[9][2]  ( .A(n15578), .EN(n15579), .Y(\regZ[9][2] ) );
  TBUFX1 \regZ_tri[9][3]  ( .A(n15580), .EN(n15581), .Y(\regZ[9][3] ) );
  TBUFX1 \regZ_tri[9][4]  ( .A(n15582), .EN(n15583), .Y(\regZ[9][4] ) );
  TBUFX1 \regZ_tri[9][5]  ( .A(n15584), .EN(n15585), .Y(\regZ[9][5] ) );
  TBUFX1 \regZ_tri[9][6]  ( .A(n15586), .EN(n15587), .Y(\regZ[9][6] ) );
  TBUFX1 \regZ_tri[9][7]  ( .A(n15588), .EN(n15589), .Y(\regZ[9][7] ) );
  TBUFX1 \regZ_tri[8][0]  ( .A(n15558), .EN(n15559), .Y(\regZ[8][0] ) );
  TBUFX1 \regZ_tri[8][1]  ( .A(n15560), .EN(n15561), .Y(\regZ[8][1] ) );
  TBUFX1 \regZ_tri[8][2]  ( .A(n15562), .EN(n15563), .Y(\regZ[8][2] ) );
  TBUFX1 \regZ_tri[8][3]  ( .A(n15564), .EN(n15565), .Y(\regZ[8][3] ) );
  TBUFX1 \regZ_tri[8][4]  ( .A(n15566), .EN(n15567), .Y(\regZ[8][4] ) );
  TBUFX1 \regZ_tri[8][5]  ( .A(n15568), .EN(n15569), .Y(\regZ[8][5] ) );
  TBUFX1 \regZ_tri[8][6]  ( .A(n15570), .EN(n15571), .Y(\regZ[8][6] ) );
  TBUFX1 \regZ_tri[8][7]  ( .A(n15572), .EN(n15573), .Y(\regZ[8][7] ) );
  TBUFX1 \regZ_tri[7][0]  ( .A(n15542), .EN(n15543), .Y(\regZ[7][0] ) );
  TBUFX1 \regZ_tri[7][1]  ( .A(n15544), .EN(n15545), .Y(\regZ[7][1] ) );
  TBUFX1 \regZ_tri[7][2]  ( .A(n15546), .EN(n15547), .Y(\regZ[7][2] ) );
  TBUFX1 \regZ_tri[7][3]  ( .A(n15548), .EN(n15549), .Y(\regZ[7][3] ) );
  TBUFX1 \regZ_tri[7][4]  ( .A(n15550), .EN(n15551), .Y(\regZ[7][4] ) );
  TBUFX1 \regZ_tri[7][5]  ( .A(n15552), .EN(n15553), .Y(\regZ[7][5] ) );
  TBUFX1 \regZ_tri[7][6]  ( .A(n15554), .EN(n15555), .Y(\regZ[7][6] ) );
  TBUFX1 \regZ_tri[7][7]  ( .A(n15556), .EN(n15557), .Y(\regZ[7][7] ) );
  TBUFX1 \regZ_tri[6][0]  ( .A(n15526), .EN(n15527), .Y(\regZ[6][0] ) );
  TBUFX1 \regZ_tri[6][1]  ( .A(n15528), .EN(n15529), .Y(\regZ[6][1] ) );
  TBUFX1 \regZ_tri[6][2]  ( .A(n15530), .EN(n15531), .Y(\regZ[6][2] ) );
  TBUFX1 \regZ_tri[6][3]  ( .A(n15532), .EN(n15533), .Y(\regZ[6][3] ) );
  TBUFX1 \regZ_tri[6][4]  ( .A(n15534), .EN(n15535), .Y(\regZ[6][4] ) );
  TBUFX1 \regZ_tri[6][5]  ( .A(n15536), .EN(n15537), .Y(\regZ[6][5] ) );
  TBUFX1 \regZ_tri[6][6]  ( .A(n15538), .EN(n15539), .Y(\regZ[6][6] ) );
  TBUFX1 \regZ_tri[6][7]  ( .A(n15540), .EN(n15541), .Y(\regZ[6][7] ) );
  TBUFX1 \regZ_tri[5][0]  ( .A(n15510), .EN(n15511), .Y(\regZ[5][0] ) );
  TBUFX1 \regZ_tri[5][1]  ( .A(n15512), .EN(n15513), .Y(\regZ[5][1] ) );
  TBUFX1 \regZ_tri[5][2]  ( .A(n15514), .EN(n15515), .Y(\regZ[5][2] ) );
  TBUFX1 \regZ_tri[5][3]  ( .A(n15516), .EN(n15517), .Y(\regZ[5][3] ) );
  TBUFX1 \regZ_tri[5][4]  ( .A(n15518), .EN(n15519), .Y(\regZ[5][4] ) );
  TBUFX1 \regZ_tri[5][5]  ( .A(n15520), .EN(n15521), .Y(\regZ[5][5] ) );
  TBUFX1 \regZ_tri[5][6]  ( .A(n15522), .EN(n15523), .Y(\regZ[5][6] ) );
  TBUFX1 \regZ_tri[5][7]  ( .A(n15524), .EN(n15525), .Y(\regZ[5][7] ) );
  TBUFX1 \regZ_tri[4][0]  ( .A(n15494), .EN(n15495), .Y(\regZ[4][0] ) );
  TBUFX1 \regZ_tri[4][1]  ( .A(n15496), .EN(n15497), .Y(\regZ[4][1] ) );
  TBUFX1 \regZ_tri[4][2]  ( .A(n15498), .EN(n15499), .Y(\regZ[4][2] ) );
  TBUFX1 \regZ_tri[4][3]  ( .A(n15500), .EN(n15501), .Y(\regZ[4][3] ) );
  TBUFX1 \regZ_tri[4][4]  ( .A(n15502), .EN(n15503), .Y(\regZ[4][4] ) );
  TBUFX1 \regZ_tri[4][5]  ( .A(n15504), .EN(n15505), .Y(\regZ[4][5] ) );
  TBUFX1 \regZ_tri[4][6]  ( .A(n15506), .EN(n15507), .Y(\regZ[4][6] ) );
  TBUFX1 \regZ_tri[4][7]  ( .A(n15508), .EN(n15509), .Y(\regZ[4][7] ) );
  TBUFX1 \regZ_tri[3][0]  ( .A(n15478), .EN(n15479), .Y(\regZ[3][0] ) );
  TBUFX1 \regZ_tri[3][1]  ( .A(n15480), .EN(n15481), .Y(\regZ[3][1] ) );
  TBUFX1 \regZ_tri[3][2]  ( .A(n15482), .EN(n15483), .Y(\regZ[3][2] ) );
  TBUFX1 \regZ_tri[3][3]  ( .A(n15484), .EN(n15485), .Y(\regZ[3][3] ) );
  TBUFX1 \regZ_tri[3][4]  ( .A(n15486), .EN(n15487), .Y(\regZ[3][4] ) );
  TBUFX1 \regZ_tri[3][5]  ( .A(n15488), .EN(n15489), .Y(\regZ[3][5] ) );
  TBUFX1 \regZ_tri[3][6]  ( .A(n15490), .EN(n15491), .Y(\regZ[3][6] ) );
  TBUFX1 \regZ_tri[3][7]  ( .A(n15492), .EN(n15493), .Y(\regZ[3][7] ) );
  TBUFX1 \regZ_tri[2][0]  ( .A(n15829), .EN(n15828), .Y(\regZ[2][0] ) );
  TBUFX1 \regZ_tri[2][1]  ( .A(n15827), .EN(n15826), .Y(\regZ[2][1] ) );
  TBUFX1 \regZ_tri[2][2]  ( .A(n15825), .EN(n15824), .Y(\regZ[2][2] ) );
  TBUFX1 \regZ_tri[2][3]  ( .A(n15823), .EN(n15822), .Y(\regZ[2][3] ) );
  TBUFX1 \regZ_tri[2][4]  ( .A(n15821), .EN(n15820), .Y(\regZ[2][4] ) );
  TBUFX1 \regZ_tri[2][5]  ( .A(n15819), .EN(n15818), .Y(\regZ[2][5] ) );
  TBUFX1 \regZ_tri[2][6]  ( .A(n15817), .EN(n15816), .Y(\regZ[2][6] ) );
  TBUFX1 \regZ_tri[2][7]  ( .A(n15815), .EN(n15814), .Y(\regZ[2][7] ) );
  TBUFX1 \regZ_tri[1][0]  ( .A(n15845), .EN(n15844), .Y(\regZ[1][0] ) );
  TBUFX1 \regZ_tri[1][1]  ( .A(n15843), .EN(n15842), .Y(\regZ[1][1] ) );
  TBUFX1 \regZ_tri[1][2]  ( .A(n15841), .EN(n15840), .Y(\regZ[1][2] ) );
  TBUFX1 \regZ_tri[1][3]  ( .A(n15839), .EN(n15838), .Y(\regZ[1][3] ) );
  TBUFX1 \regZ_tri[1][4]  ( .A(n15837), .EN(n15836), .Y(\regZ[1][4] ) );
  TBUFX1 \regZ_tri[1][5]  ( .A(n15835), .EN(n15834), .Y(\regZ[1][5] ) );
  TBUFX1 \regZ_tri[1][6]  ( .A(n15833), .EN(n15832), .Y(\regZ[1][6] ) );
  TBUFX1 \regZ_tri[1][7]  ( .A(n15831), .EN(n15830), .Y(\regZ[1][7] ) );
  TBUFX1 \regZ_tri[0][0]  ( .A(n15411), .EN(n15412), .Y(\regZ[0][0] ) );
  TBUFX1 \regZ_tri[0][1]  ( .A(n15413), .EN(n15414), .Y(\regZ[0][1] ) );
  TBUFX1 \regZ_tri[0][2]  ( .A(n15415), .EN(n15416), .Y(\regZ[0][2] ) );
  TBUFX1 \regZ_tri[0][3]  ( .A(n15417), .EN(n15418), .Y(\regZ[0][3] ) );
  TBUFX1 \regZ_tri[0][4]  ( .A(n15426), .EN(n15425), .Y(\regZ[0][4] ) );
  TBUFX1 \regZ_tri[0][5]  ( .A(n15424), .EN(n15423), .Y(\regZ[0][5] ) );
  TBUFX1 \regZ_tri[0][6]  ( .A(n15422), .EN(n15421), .Y(\regZ[0][6] ) );
  TBUFX1 \regZ_tri[0][7]  ( .A(n15420), .EN(n15419), .Y(\regZ[0][7] ) );
  CannyEdge_DW01_addsub_1 add_0_root_add_205_8 ( .A({N2416, N2415, N2414, 
        N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, 
        N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, 
        N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385}), .B({
        N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, 
        N2470, N2469, N2468, N2467, N2466, N2465, N2464, N1912, N1911, N1910, 
        N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, 
        N1899, N1898}), .CI(1'b0), .ADD_SUB(1'b0), .SUM({N2544, N2543, N2542, 
        N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, 
        N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, 
        N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513}) );
  CannyEdge_DW01_addsub_3 add_0_root_add_160_24 ( .A({N2002, N2001, N2000, 
        N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, 
        N1989, N1988}), .B({N2032, N2031, N2030, N2029, N2028, N2027, N2026, 
        N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N2055, N2054, N2053, N2052, N2051, N2050, N2049, 
        N2048, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  CannyEdge_DW01_addsub_4 add_1_root_add_160_24 ( .A({N1942, N1941, N1940, 
        N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, 
        N1929, N1928}), .B({N1972, N1971, N1970, N1969, N1968, N1967, N1966, 
        N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N2032, N2031, N2030, N2029, N2028, N2027, N2026, 
        N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018}) );
  CannyEdge_DW01_add_0 add_3_root_add_160_24 ( .A({N1822, N1821, N1820, N1819, 
        N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, 
        1'b0}), .B({N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, 
        N1844, N1843, N1842, N1841, N1840, N1839, N1838}), .CI(1'b0), .SUM({
        N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, 
        N1962, N1961, N1960, N1959, N1958}) );
  CannyEdge_DW01_add_1 add_7_root_add_160_24 ( .A({N1582, N1581, N1580, N1579, 
        N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, 
        N1568}), .B({N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, 
        N1604, N1603, N1602, N1601, N1600, N1599, N1598}), .CI(1'b0), .SUM({
        N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, 
        N1842, N1841, N1840, N1839, N1838}) );
  CannyEdge_DW01_add_2 add_15_root_add_160_24 ( .A({1'b0, N1806, N1805, N1804, 
        N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, 
        N1793}), .B({1'b0, N1836, N1835, N1834, N1833, N1832, N1831, N1830, 
        N1829, N1828, N1827, N1826, N1825, N1824, 1'b0}), .CI(1'b0), .SUM({
        N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, 
        N1602, N1601, N1600, N1599, N1598}) );
  CannyEdge_DW01_add_4 add_8_root_add_160_24 ( .A({N1522, N1521, N1520, N1519, 
        N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, 
        1'b0}), .B({N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, 
        N1544, N1543, N1542, N1541, N1540, N1539, 1'b0}), .CI(1'b0), .SUM({
        N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, 
        N1812, N1811, N1810, N1809, SYNOPSYS_UNCONNECTED__7}) );
  CannyEdge_DW01_add_7 add_4_root_add_160_24 ( .A({N1762, N1761, N1760, N1759, 
        N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, 
        N1748}), .B({N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, 
        N1784, N1783, N1782, N1781, N1780, N1779, N1778}), .CI(1'b0), .SUM({
        N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, 
        N1932, N1931, N1930, N1929, N1928}) );
  CannyEdge_DW01_add_8 add_9_root_add_160_24 ( .A({N1462, N1461, N1460, N1459, 
        N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, 
        N1448}), .B({N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, 
        N1484, N1483, N1482, N1481, N1480, N1479, N1478}), .CI(1'b0), .SUM({
        N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, 
        N1782, N1781, N1780, N1779, N1778}) );
  CannyEdge_DW01_add_9 add_19_root_add_160_24 ( .A({1'b0, N1566, N1565, N1564, 
        N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, 
        N1553}), .B({1'b0, N1596, N1595, N1594, N1593, N1592, N1591, N1590, 
        N1589, N1588, N1587, N1586, N1585, N1584, N1583}), .CI(1'b0), .SUM({
        N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, 
        N1482, N1481, N1480, N1479, N1478}) );
  CannyEdge_DW01_add_10 add_10_root_add_160_24 ( .A({N1402, N1401, N1400, 
        N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, 
        N1389, N1388}), .B({N2186, N2185, N2184, N2183, N2182, N2181, N2180, 
        N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172}), .CI(1'b0), 
        .SUM({N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, 
        N1753, N1752, N1751, N1750, N1749, N1748}) );
  CannyEdge_DW01_add_11 add_2_root_add_160_24 ( .A({N1882, N1881, N1880, N1879, 
        N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, 
        N1868}), .B({N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, 
        N1904, N1903, N1902, N1901, N1900, N1899, N1898}), .CI(1'b0), .SUM({
        N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, 
        N1992, N1991, N1990, N1989, N1988}) );
  CannyEdge_DW01_add_12 r1417 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U76/Z_14 , \U3/U76/Z_13 , \U3/U76/Z_12 , \U3/U76/Z_11 , 
        \U3/U76/Z_10 , n15329, n15330, n15331, n15356, n15357, n15358, n15359, 
        n15360, n15361, n15362}), .B({\U3/U77/Z_31 , \U3/U77/Z_30 , 
        \U3/U77/Z_29 , \U3/U77/Z_28 , \U3/U77/Z_27 , \U3/U77/Z_26 , 
        \U3/U77/Z_25 , \U3/U77/Z_24 , \U3/U77/Z_23 , \U3/U77/Z_22 , 
        \U3/U77/Z_21 , \U3/U77/Z_20 , \U3/U77/Z_19 , \U3/U77/Z_18 , 
        \U3/U77/Z_17 , \U3/U77/Z_16 , \U3/U77/Z_15 , N1732, N1731, N1730, 
        N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, 
        N1719, N1718}), .CI(1'b0), .SUM({N2480, N2479, N2478, N2477, N2476, 
        N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, 
        N2465, N2464, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, 
        N1904, N1903, N1902, N1901, N1900, N1899, N1898}) );
  CannyEdge_DW01_add_13 add_4_root_add_205_8 ( .A({1'b0, 1'b0, \regX[0][7] , 
        \regX[0][6] , \regX[0][5] , \regX[0][4] , \regX[0][3] , \regX[0][2] , 
        \regX[0][1] , \regX[0][0] }), .B({1'b0, \regX[1][7] , \regX[1][6] , 
        \regX[1][5] , \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] , 
        \regX[1][0] , 1'b0}), .CI(1'b0), .SUM({N2341, N2340, N2339, N2338, 
        N2337, N2336, N2335, N2334, N2333, N2332}) );
  CannyEdge_DW01_add_14 r1263 ( .A({\U3/U74/Z_31 , \U3/U74/Z_30 , 
        \U3/U74/Z_29 , \U3/U74/Z_28 , \U3/U74/Z_27 , \U3/U74/Z_26 , 
        \U3/U74/Z_25 , \U3/U74/Z_24 , \U3/U74/Z_23 , \U3/U74/Z_22 , 
        \U3/U74/Z_21 , \U3/U74/Z_20 , \U3/U74/Z_19 , \U3/U74/Z_18 , 
        \U3/U74/Z_17 , \U3/U74/Z_16 , \U3/U74/Z_15 , N2250, N2249, N2248, 
        N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, 
        N2237, N2236}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \U3/U75/Z_14 , 
        \U3/U75/Z_13 , \U3/U75/Z_12 , \U3/U75/Z_11 , \U3/U75/Z_10 , 
        \U3/U75/Z_9 , \U3/U75/Z_8 , \U3/U75/Z_7 , \U3/U75/Z_6 , \U3/U75/Z_5 , 
        \U3/U75/Z_4 , \U3/U75/Z_3 , \U3/U75/Z_2 , \U3/U75/Z_1 , \U3/U75/Z_0 }), 
        .CI(1'b0), .SUM({\U3/U77/DATA2_31 , \U3/U77/DATA2_30 , 
        \U3/U77/DATA2_29 , \U3/U77/DATA2_28 , \U3/U77/DATA2_27 , 
        \U3/U77/DATA2_26 , \U3/U77/DATA2_25 , \U3/U77/DATA2_24 , 
        \U3/U77/DATA2_23 , \U3/U77/DATA2_22 , \U3/U77/DATA2_21 , 
        \U3/U77/DATA2_20 , \U3/U77/DATA2_19 , \U3/U77/DATA2_18 , 
        \U3/U77/DATA2_17 , \U3/U77/DATA2_16 , \U3/U77/DATA2_15 , N1732, N1731, 
        N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, 
        N1720, N1719, N1718}) );
  CannyEdge_DW01_add_15 r1259 ( .A({\U3/U72/Z_31 , \U3/U72/Z_30 , 
        \U3/U72/Z_29 , \U3/U72/Z_28 , \U3/U72/Z_27 , \U3/U72/Z_26 , 
        \U3/U72/Z_25 , \U3/U72/Z_24 , \U3/U72/Z_23 , \U3/U72/Z_22 , 
        \U3/U72/Z_21 , \U3/U72/Z_20 , \U3/U72/Z_19 , \U3/U72/Z_18 , 
        \U3/U72/Z_17 , \U3/U72/Z_16 , \U3/U72/Z_15 , N2823, N2822, N2821, 
        N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, 
        N2810, N2417}), .B({\U3/U73/Z_31 , \U3/U73/Z_30 , \U3/U73/Z_29 , 
        \U3/U73/Z_28 , \U3/U73/Z_27 , \U3/U73/Z_26 , \U3/U73/Z_25 , 
        \U3/U73/Z_24 , \U3/U73/Z_23 , \U3/U73/Z_22 , \U3/U73/Z_21 , 
        \U3/U73/Z_20 , \U3/U73/Z_19 , \U3/U73/Z_18 , \U3/U73/Z_17 , 
        \U3/U73/Z_16 , \U3/U73/Z_15 , N2894, N2893, N2892, N2891, N2890, N2889, 
        N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2481}), .CI(
        1'b0), .SUM({N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, 
        N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, 
        N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, 
        N2388, N2387, N2386, N2385}) );
  CannyEdge_DW01_add_16 add_6_root_add_160_24 ( .A({N1642, N1641, N1640, N1639, 
        N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, 
        N1628}), .B({N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, 
        N1664, N1663, N1662, N1661, N1660, N1659, N1658}), .CI(1'b0), .SUM({
        N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, 
        N1872, N1871, N1870, N1869, N1868}) );
  CannyEdge_DW01_add_17 add_13_root_add_160_24 ( .A({N1927, N1926, N1925, 
        N1924, N1923, N1922, N1921, N1920, N1919, N1918, N3093, N3092, N3091, 
        N3090, N3089}), .B({N1957, N1956, N1955, N1954, N1953, N1952, N1951, 
        N1950, N1949, N3194, N3193, N3192, N3191, N3190, N3189}), .CI(1'b0), 
        .SUM({N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, 
        N1663, N1662, N1661, N1660, N1659, N1658}) );
  CannyEdge_DW01_add_18 add_14_root_add_160_24 ( .A({N1867, N1866, N1865, 
        N1864, N1863, N1862, N1861, N1860, N1859, N1858, N3343, N3342, N3341, 
        N3340, N3359}), .B({1'b0, N1896, N1895, N1894, N1893, N1892, N1891, 
        N1890, N1889, N976, N975, N974, N973, N972, N971}), .CI(1'b0), .SUM({
        N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, 
        N1632, N1631, N1630, N1629, N1628}) );
  CannyEdge_DW01_addsub_5 add_20_root_add_160_24 ( .A({1'b0, N1506, N1505, 
        N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, 
        N1494, N1493}), .B({1'b0, N1536, N1535, N1534, N1533, N1532, N1531, 
        N1530, N1529, N1528, N1527, N1526, N1525, N1524, 1'b0}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N1462, N1461, N1460, N1459, N1458, N1457, N1456, 
        N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448}) );
  CannyEdge_DW01_addsub_7 r1802 ( .A({\U3/U78/Z_31 , \U3/U78/Z_30 , 
        \U3/U78/Z_29 , \U3/U78/Z_28 , \U3/U78/Z_27 , \U3/U78/Z_26 , 
        \U3/U78/Z_25 , \U3/U78/Z_24 , \U3/U78/Z_23 , \U3/U78/Z_22 , 
        \U3/U78/Z_21 , \U3/U78/Z_20 , \U3/U78/Z_19 , \U3/U78/Z_18 , 
        \U3/U78/Z_17 , \U3/U78/Z_16 , \U3/U78/Z_15 , \U3/U78/Z_14 , 
        \U3/U78/Z_13 , \U3/U78/Z_12 , \U3/U78/Z_11 , \U3/U78/Z_10 , 
        \U3/U78/Z_9 , \U3/U78/Z_8 , \U3/U78/Z_7 , \U3/U78/Z_6 , \U3/U78/Z_5 , 
        \U3/U78/Z_4 , \U3/U78/Z_3 , \U3/U78/Z_2 , \U3/U78/Z_1 , \U3/U78/Z_0 }), 
        .B({\U3/U79/Z_31 , \U3/U79/Z_30 , \U3/U79/Z_29 , \U3/U79/Z_28 , 
        \U3/U79/Z_27 , \U3/U79/Z_26 , \U3/U79/Z_25 , \U3/U79/Z_24 , 
        \U3/U79/Z_23 , \U3/U79/Z_22 , \U3/U79/Z_21 , \U3/U79/Z_20 , 
        \U3/U79/Z_19 , \U3/U79/Z_18 , \U3/U79/Z_17 , \U3/U79/Z_16 , 
        \U3/U79/Z_15 , \U3/U79/Z_14 , \U3/U79/Z_13 , \U3/U79/Z_12 , 
        \U3/U79/Z_11 , \U3/U79/Z_10 , \U3/U79/Z_9 , \U3/U79/Z_8 , \U3/U79/Z_7 , 
        \U3/U79/Z_6 , \U3/U79/Z_5 , \U3/U79/Z_4 , \U3/U79/Z_3 , \U3/U79/Z_2 , 
        \U3/U79/Z_1 , \U3/U79/Z_0 }), .CI(1'b0), .ADD_SUB(n12475), .SUM({N2331, 
        N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, 
        N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, 
        N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, 
        N2300}) );
  CannyEdge_DW01_add_19 add_1_root_add_202_8 ( .A({N2139, N2138, N2137, N2136, 
        N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, 
        N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, 
        N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108}), .B({N2203, 
        N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, 
        N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, 
        N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, 
        N2172}), .CI(1'b0), .SUM({N2299, N2298, N2297, N2296, N2295, N2294, 
        N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, 
        N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, 
        N2273, N2272, N2271, N2270, N2269, N2268}) );
  CannyEdge_DW01_add_20 r1223 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \U3/U70/Z_8 , \U3/U70/Z_7 , \U3/U70/Z_6 , 
        \U3/U70/Z_5 , \U3/U70/Z_4 , \U3/U70/Z_3 , \U3/U70/Z_2 , \U3/U70/Z_1 , 
        \U3/U70/Z_0 }), .B({\U3/U71/Z_31 , \U3/U71/Z_30 , \U3/U71/Z_29 , 
        \U3/U71/Z_28 , \U3/U71/Z_27 , \U3/U71/Z_26 , \U3/U71/Z_25 , 
        \U3/U71/Z_24 , \U3/U71/Z_23 , \U3/U71/Z_22 , \U3/U71/Z_21 , 
        \U3/U71/Z_20 , \U3/U71/Z_19 , \U3/U71/Z_18 , \U3/U71/Z_17 , 
        \U3/U71/Z_16 , \U3/U71/Z_15 , N2154, N2153, N2152, N2151, N2150, N2149, 
        N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140}), .CI(
        1'b0), .SUM({N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, 
        N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, 
        N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, 
        N2175, N2174, N2173, N2172}) );
  CannyEdge_DW01_add_21 r1814 ( .A({\U3/U68/Z_31 , \U3/U68/Z_30 , 
        \U3/U68/Z_29 , \U3/U68/Z_28 , \U3/U68/Z_27 , \U3/U68/Z_26 , 
        \U3/U68/Z_25 , \U3/U68/Z_24 , \U3/U68/Z_23 , \U3/U68/Z_22 , 
        \U3/U68/Z_21 , \U3/U68/Z_20 , \U3/U68/Z_19 , \U3/U68/Z_18 , 
        \U3/U68/Z_17 , \U3/U68/Z_16 , \U3/U68/Z_15 , N2090, N2089, N2088, 
        N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, 
        N2077, N2076}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U69/Z_13 , \U3/U69/Z_12 , \U3/U69/Z_11 , \U3/U69/Z_10 , 
        \U3/U69/Z_9 , \U3/U69/Z_8 , \U3/U69/Z_7 , \U3/U69/Z_6 , \U3/U69/Z_5 , 
        \U3/U69/Z_4 , \U3/U69/Z_3 , \U3/U69/Z_2 , \U3/U69/Z_1 , \U3/U69/Z_0 }), 
        .CI(1'b0), .SUM({N2139, N2138, N2137, N2136, N2135, N2134, N2133, 
        N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, 
        N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, 
        N2112, N2111, N2110, N2109, N2108}) );
  CannyEdge_DW01_addsub_9 r1201 ( .A({\U3/U100/Z_6 , n15326, \U3/U100/Z_4 , 
        \U3/U100/Z_3 , \U3/U100/Z_2 , \U3/U100/Z_1 , \U3/U100/Z_0 }), .B({
        \U3/U101/Z_6 , \U3/U101/Z_6 , \U3/U101/Z_6 , \U3/U101/Z_3 , 
        \U3/U101/Z_2 , \U3/U101/Z_1 , \U3/U101/Z_0 }), .CI(1'b0), .ADD_SUB(
        1'b0), .SUM({N983, N982, N981, N980, N979, N978, N977}) );
  CannyEdge_DW01_addsub_11 r1337 ( .A({\U3/U134/Z_10 , \U3/U134/Z_9 , 
        \U3/U134/Z_8 , \U3/U134/Z_7 , \U3/U134/Z_6 , \U3/U134/Z_5 , 
        \U3/U134/Z_4 , \U3/U134/Z_3 , \U3/U134/Z_2 , \U3/U134/Z_1 , 
        \U3/U134/Z_0 }), .B({n12449, n12450, n12451, n12452, n12453, n12454, 
        n12455, n12456, n12457, n12458, n12459}), .CI(1'b0), .ADD_SUB(
        \U3/U136/Z_0 ), .SUM({N2576, N2575, N2574, N2573, N2572, N2571, N2570, 
        N2569, SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  CannyEdge_DW01_addsub_12 r1343 ( .A(Gx[10:0]), .B(Gy[10:0]), .CI(1'b0), 
        .ADD_SUB(n8303), .SUM({N2568, N2567, N2566, N2565, N2564, N2563, N2562, 
        N2561, N2560, N2559, N2558}) );
  CannyEdge_DW01_cmp2_0 lte_289 ( .A(fGy), .B({N2840, N2840, N2839, N2838, 
        N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, 
        N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, 
        N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810}), .LEQ(1'b1), 
        .TC(1'b1), .LT_LE(N2841) );
  CannyEdge_DW01_cmp2_1 gt_274 ( .A({N2911, N2911, N2910, N2909, N2908, N2907, 
        N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, 
        N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, 
        N2886, N2885, N2884, N2883, N2882, N2881}), .B(fGy), .LEQ(1'b0), .TC(
        1'b1), .LT_LE(N2945) );
  CannyEdge_DW01_cmp2_2 gt_292 ( .A({N2840, N2840, N2839, N2838, N2837, N2836, 
        N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, 
        N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, 
        N2815, N2814, N2813, N2812, N2811, N2810}), .B(fGy), .LEQ(1'b0), .TC(
        1'b1), .LT_LE(N2874) );
  CannyEdge_DW02_mult_0 mult_160_18 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[17][7] , \regX[17][6] , \regX[17][5] , 
        \regX[17][4] , \regX[17][3] , \regX[17][2] , \regX[17][1] , 
        \regX[17][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, N1836, N1835, N1834, N1833, N1832, N1831, 
        N1830, N1829, N1828, N1827, N1826, N1825, N1824, 
        SYNOPSYS_UNCONNECTED__13}) );
  CannyEdge_DW02_mult_1 mult_160_17 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[16][7] , \regX[16][6] , \regX[16][5] , 
        \regX[16][4] , \regX[16][3] , \regX[16][2] , \regX[16][1] , 
        \regX[16][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N1806, N1805, N1804, N1803, N1802, N1801, 
        N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793}) );
  CannyEdge_DW02_mult_2 mult_160_16 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[15][7] , \regX[15][6] , \regX[15][5] , 
        \regX[15][4] , \regX[15][3] , \regX[15][2] , \regX[15][1] , 
        \regX[15][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, N1776, N1775, N1774, N1773, N1772, N1771, 
        N1770, N1769, N1768, N1767, N1766, N1765, N1569, N1568}) );
  CannyEdge_DW02_mult_4 mult_160_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[13][7] , \regX[13][6] , \regX[13][5] , 
        \regX[13][4] , \regX[13][3] , \regX[13][2] , \regX[13][1] , 
        \regX[13][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, N1716, N1715, N1714, N1713, N1712, N1711, 
        N1710, N1709, N1708, N1707, N1541, N1540, N1539, 
        SYNOPSYS_UNCONNECTED__20}) );
  CannyEdge_DW02_mult_6 mult_160_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[11][7] , \regX[11][6] , \regX[11][5] , 
        \regX[11][4] , \regX[11][3] , \regX[11][2] , \regX[11][1] , 
        \regX[11][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, N1656, N1655, N1654, N1653, N1652, N1651, 
        N1650, N1649, N1648, N1647, N1646, N1645, N1509, 
        SYNOPSYS_UNCONNECTED__23}) );
  CannyEdge_DW02_mult_8 mult_160_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[9][7] , \regX[9][6] , \regX[9][5] , 
        \regX[9][4] , \regX[9][3] , \regX[9][2] , \regX[9][1] , \regX[9][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, N1596, N1595, N1594, N1593, N1592, N1591, 
        N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583}) );
  CannyEdge_DW02_mult_9 mult_160_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[8][7] , \regX[8][6] , \regX[8][5] , 
        \regX[8][4] , \regX[8][3] , \regX[8][2] , \regX[8][1] , \regX[8][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N1566, N1565, N1564, N1563, N1562, N1561, 
        N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553}) );
  CannyEdge_DW02_mult_10 mult_160_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[7][7] , \regX[7][6] , \regX[7][5] , 
        \regX[7][4] , \regX[7][3] , \regX[7][2] , \regX[7][1] , \regX[7][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, N1536, N1535, N1534, N1533, N1532, N1531, 
        N1530, N1529, N1528, N1527, N1526, N1525, N1524, 
        SYNOPSYS_UNCONNECTED__30}) );
  CannyEdge_DW02_mult_11 r1229 ( .A({n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12476, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, \U3/U67/Z_1 , 
        n15370}), .B({\regX[5][7] , \regX[5][6] , \regX[5][5] , \regX[5][4] , 
        \regX[5][3] , \regX[5][2] , \regX[5][1] , \regX[5][0] }), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, N2171, N2170, 
        N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, 
        N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, 
        N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140})
         );
  CannyEdge_DW02_mult_14 mult_160_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[1][7] , \regX[1][6] , \regX[1][5] , 
        \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] , \regX[1][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, N1356, N1355, N1354, N1353, N1352, N1351, 
        N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343}) );
  CannyEdge_DW02_mult_15 r1211 ( .A({n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12476, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, 
        \U3/U67/Z_1 }), .B({\regX[0][7] , \regX[0][6] , \regX[0][5] , 
        \regX[0][4] , \regX[0][3] , \regX[0][2] , \regX[0][1] , \regX[0][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, N2107, N2106, N2105, N2104, N2103, N2102, 
        N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, 
        N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, 
        N2081, N2080, N2079, N2078, N2077, N2076}) );
  CannyEdge_DW02_mult_16 r1207 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n5396, 
        n5397, n5398}), .B({\U3/U63/Z_7 , \U3/U63/Z_6 , \U3/U63/Z_5 , 
        \U3/U63/Z_4 , \U3/U63/Z_3 , \U3/U63/Z_2 , \U3/U63/Z_1 , \U3/U63/Z_0 }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, N1896, N1895, N1894, N1893, N1892, N1891, 
        N1890, N1889, N976, N975, N974, N973, N972, N971}) );
  CannyEdge_DW02_mult_17 r1075 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n15325, 
        n15370, \U3/U124/Z_0 }), .B({\U3/U125/Z_7 , \U3/U125/Z_6 , 
        \U3/U125/Z_5 , \U3/U125/Z_4 , \U3/U125/Z_3 , \U3/U125/Z_2 , 
        \U3/U125/Z_1 , \U3/U125/Z_0 }), .TC(n15325), .PRODUCT({
        SYNOPSYS_UNCONNECTED__51, N1417, N1416, N1415, N1414, N1413, N1412, 
        N1411, N1410, N1409, N1408, N3443, N3442, N3441, N1389, N1388}) );
  CannyEdge_DW02_mult_18 r1062 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n15327, 
        n15370, \U3/U97/Z_0 }), .B({\U3/U98/Z_7 , \U3/U98/Z_6 , \U3/U98/Z_5 , 
        \U3/U98/Z_4 , \U3/U98/Z_3 , \U3/U98/Z_2 , \U3/U98/Z_1 , \U3/U98/Z_0 }), 
        .TC(n15327), .PRODUCT({SYNOPSYS_UNCONNECTED__52, N1957, N1956, N1955, 
        N1954, N1953, N1952, N1951, N1950, N1949, N3194, N3193, N3192, N3191, 
        N3190, N3189}) );
  CannyEdge_DW01_cmp2_3 r1050 ( .A({n15334, n15335, n15336, n15337, n15338, 
        n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, 
        n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15332, 
        n15333, \U3/U121/Z_7 , \U3/U121/Z_6 , \U3/U121/Z_5 , \U3/U121/Z_4 , 
        \U3/U121/Z_3 , \U3/U121/Z_2 , \U3/U121/Z_1 , \U3/U121/Z_0 }), .B({1'b0, 
        1'b0, \U3/U122/Z_29 , \U3/U122/Z_28 , \U3/U122/Z_27 , \U3/U122/Z_26 , 
        \U3/U122/Z_25 , \U3/U122/Z_24 , \U3/U122/Z_23 , \U3/U122/Z_22 , 
        \U3/U122/Z_21 , \U3/U122/Z_20 , \U3/U122/Z_19 , \U3/U122/Z_18 , 
        \U3/U122/Z_17 , \U3/U122/Z_16 , \U3/U122/Z_15 , \U3/U122/Z_14 , 
        \U3/U122/Z_13 , \U3/U122/Z_12 , \U3/U122/Z_11 , \U3/U122/Z_10 , 
        \U3/U122/Z_9 , \U3/U122/Z_8 , \U3/U122/Z_7 , \U3/U122/Z_6 , 
        \U3/U122/Z_5 , \U3/U122/Z_4 , \U3/U122/Z_3 , \U3/U122/Z_2 , 
        \U3/U122/Z_1 , \U3/U122/Z_0 }), .LEQ(1'b1), .TC(n12466), .GE_GT(N2880)
         );
  CannyEdge_DW02_mult_19 r1047 ( .A({\U3/U84/Z_7 , \U3/U84/Z_6 , \U3/U84/Z_5 , 
        \U3/U84/Z_4 , \U3/U84/Z_3 , \U3/U84/Z_2 , \U3/U84/Z_1 , \U3/U84/Z_0 }), 
        .B({\U3/U85/Z_31 , \U3/U85/Z_30 , \U3/U85/Z_29 , \U3/U85/Z_28 , 
        \U3/U85/Z_27 , \U3/U85/Z_26 , \U3/U85/Z_25 , \U3/U85/Z_24 , 
        \U3/U85/Z_23 , \U3/U85/Z_22 , \U3/U85/Z_21 , \U3/U85/Z_20 , 
        \U3/U85/Z_19 , \U3/U85/Z_18 , \U3/U85/Z_17 , \U3/U85/Z_16 , 
        \U3/U85/Z_15 , \U3/U85/Z_14 , \U3/U85/Z_13 , \U3/U85/Z_12 , 
        \U3/U85/Z_11 , \U3/U85/Z_10 , \U3/U85/Z_9 , \U3/U85/Z_8 , \U3/U85/Z_7 , 
        \U3/U85/Z_6 , \U3/U85/Z_5 , \U3/U85/Z_4 , \U3/U85/Z_3 , \U3/U85/Z_2 , 
        \U3/U85/Z_1 , \U3/U85/Z_0 }), .TC(n15377), .PRODUCT({
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, N2840, N2839, 
        N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, 
        N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, 
        N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2417})
         );
  CannyEdge_DW01_cmp2_4 r1033 ( .A({\U3/U93/Z_31 , \U3/U93/Z_30 , 
        \U3/U93/Z_29 , \U3/U93/Z_28 , \U3/U93/Z_27 , \U3/U93/Z_26 , 
        \U3/U93/Z_25 , \U3/U93/Z_24 , \U3/U93/Z_23 , \U3/U93/Z_22 , 
        \U3/U93/Z_21 , \U3/U93/Z_20 , \U3/U93/Z_19 , \U3/U93/Z_18 , 
        \U3/U93/Z_17 , \U3/U93/Z_16 , \U3/U93/Z_15 , \U3/U93/Z_14 , 
        \U3/U93/Z_13 , \U3/U93/Z_12 , \U3/U93/Z_11 , \U3/U93/Z_10 , 
        \U3/U93/Z_9 , \U3/U93/Z_8 , \U3/U93/Z_7 , \U3/U93/Z_6 , \U3/U93/Z_5 , 
        \U3/U93/Z_4 , \U3/U93/Z_3 , \U3/U93/Z_2 , \U3/U93/Z_1 , \U3/U93/Z_0 }), 
        .B({\U3/U94/Z_31 , \U3/U94/Z_31 , \U3/U94/Z_29 , \U3/U94/Z_28 , 
        \U3/U94/Z_27 , \U3/U94/Z_26 , \U3/U94/Z_25 , \U3/U94/Z_24 , 
        \U3/U94/Z_23 , \U3/U94/Z_22 , \U3/U94/Z_21 , \U3/U94/Z_20 , 
        \U3/U94/Z_19 , \U3/U94/Z_18 , \U3/U94/Z_17 , \U3/U94/Z_16 , 
        \U3/U94/Z_15 , \U3/U94/Z_14 , \U3/U94/Z_13 , \U3/U94/Z_12 , 
        \U3/U94/Z_11 , \U3/U94/Z_10 , \U3/U94/Z_9 , \U3/U94/Z_8 , \U3/U94/Z_7 , 
        \U3/U94/Z_6 , \U3/U94/Z_5 , \U3/U94/Z_4 , \U3/U94/Z_3 , \U3/U94/Z_2 , 
        \U3/U94/Z_1 , \U3/U94/Z_0 }), .LEQ(\U3/U95/Z_0 ), .TC(\U3/U96/Z_0 ), 
        .GE_GT(N2549) );
  CannyEdge_DW02_mult_20 r1051 ( .A({\U3/U87/Z_7 , \U3/U87/Z_6 , \U3/U87/Z_5 , 
        \U3/U87/Z_4 , \U3/U87/Z_3 , \U3/U87/Z_2 , \U3/U87/Z_1 , \U3/U87/Z_0 }), 
        .B({n12476, \U3/U88/Z_30 , \U3/U88/Z_29 , \U3/U88/Z_28 , \U3/U88/Z_27 , 
        \U3/U88/Z_26 , \U3/U88/Z_25 , \U3/U88/Z_24 , \U3/U88/Z_23 , 
        \U3/U88/Z_22 , \U3/U88/Z_21 , \U3/U88/Z_20 , \U3/U88/Z_19 , 
        \U3/U88/Z_18 , \U3/U88/Z_17 , \U3/U88/Z_16 , \U3/U88/Z_15 , 
        \U3/U88/Z_14 , \U3/U88/Z_13 , \U3/U88/Z_12 , \U3/U88/Z_11 , 
        \U3/U88/Z_10 , \U3/U88/Z_9 , \U3/U88/Z_8 , \U3/U88/Z_7 , \U3/U88/Z_6 , 
        \U3/U88/Z_5 , \U3/U88/Z_4 , \U3/U88/Z_3 , \U3/U88/Z_2 , \U3/U88/Z_1 , 
        \U3/U88/Z_0 }), .TC(n12466), .PRODUCT({SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, N2911, N2910, N2909, N2908, N2907, N2906, 
        N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, 
        N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, 
        N2885, N2884, N2883, N2882, N2881, N2481}) );
  CannyEdge_DW02_mult_21 mult_160_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[6][7] , \regX[6][6] , \regX[6][5] , 
        \regX[6][4] , \regX[6][3] , \regX[6][2] , \regX[6][1] , \regX[6][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, N1506, N1505, N1504, N1503, N1502, N1501, 
        N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493}) );
  CannyEdge_DW01_cmp2_5 r169 ( .A({\U3/U118/Z_31 , \U3/U118/Z_30 , 
        \U3/U118/Z_29 , \U3/U118/Z_28 , \U3/U118/Z_27 , \U3/U118/Z_26 , 
        \U3/U118/Z_25 , \U3/U118/Z_24 , \U3/U118/Z_23 , \U3/U118/Z_22 , 
        \U3/U118/Z_21 , \U3/U118/Z_20 , \U3/U118/Z_19 , \U3/U118/Z_18 , 
        \U3/U118/Z_17 , \U3/U118/Z_16 , \U3/U118/Z_15 , \U3/U118/Z_14 , 
        \U3/U118/Z_13 , \U3/U118/Z_12 , \U3/U118/Z_11 , \U3/U118/Z_10 , 
        \U3/U118/Z_9 , \U3/U118/Z_8 , \U3/U118/Z_7 , \U3/U118/Z_6 , 
        \U3/U118/Z_5 , \U3/U118/Z_4 , \U3/U118/Z_3 , \U3/U118/Z_2 , 
        \U3/U118/Z_1 , \U3/U118/Z_0 }), .B({\U3/U119/Z_31 , \U3/U119/Z_31 , 
        \U3/U119/Z_29 , \U3/U119/Z_28 , \U3/U119/Z_27 , \U3/U119/Z_26 , 
        \U3/U119/Z_25 , \U3/U119/Z_24 , \U3/U119/Z_23 , \U3/U119/Z_22 , 
        \U3/U119/Z_21 , \U3/U119/Z_20 , \U3/U119/Z_19 , \U3/U119/Z_18 , 
        \U3/U119/Z_17 , \U3/U119/Z_16 , \U3/U119/Z_15 , \U3/U119/Z_14 , 
        \U3/U119/Z_13 , \U3/U119/Z_12 , \U3/U119/Z_11 , \U3/U119/Z_10 , 
        \U3/U119/Z_9 , \U3/U119/Z_8 , \U3/U119/Z_7 , \U3/U119/Z_6 , 
        \U3/U119/Z_5 , \U3/U119/Z_4 , \U3/U119/Z_3 , \U3/U119/Z_2 , 
        \U3/U119/Z_1 , \U3/U119/Z_0 }), .LEQ(1'b1), .TC(n15377), .LT_LE(N2777)
         );
  CannyEdge_DW02_mult_22 r1055 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n15369, 
        1'b0, \U3/U90/Z_0 }), .B({\U3/U91/Z_7 , \U3/U91/Z_6 , \U3/U91/Z_5 , 
        \U3/U91/Z_4 , \U3/U91/Z_3 , \U3/U91/Z_2 , \U3/U91/Z_1 , \U3/U91/Z_0 }), 
        .TC(n15369), .PRODUCT({SYNOPSYS_UNCONNECTED__71, N1927, N1926, N1925, 
        N1924, N1923, N1922, N1921, N1920, N1919, N1918, N3093, N3092, N3091, 
        N3090, N3089}) );
  CannyEdge_DW02_mult_23 r1068 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U109/Z_2 , n15370, \U3/U109/Z_2 }), .B({\U3/U110/Z_7 , 
        \U3/U110/Z_6 , \U3/U110/Z_5 , \U3/U110/Z_4 , \U3/U110/Z_3 , 
        \U3/U110/Z_2 , \U3/U110/Z_1 , n5409}), .TC(n15328), .PRODUCT({
        SYNOPSYS_UNCONNECTED__72, N1867, N1866, N1865, N1864, N1863, N1862, 
        N1861, N1860, N1859, N1858, N3343, N3342, N3341, N3340, N3359}) );
  CannyEdge_DW01_cmp2_6 r1377 ( .A({\U3/U119/Z_31 , \U3/U119/Z_31 , 
        \U3/U119/Z_29 , \U3/U119/Z_28 , \U3/U119/Z_27 , \U3/U119/Z_26 , 
        \U3/U119/Z_25 , \U3/U119/Z_24 , \U3/U119/Z_23 , \U3/U119/Z_22 , 
        \U3/U119/Z_21 , \U3/U119/Z_20 , \U3/U119/Z_19 , \U3/U119/Z_18 , 
        \U3/U119/Z_17 , \U3/U119/Z_16 , \U3/U119/Z_15 , \U3/U119/Z_14 , 
        \U3/U119/Z_13 , \U3/U119/Z_12 , \U3/U119/Z_11 , \U3/U119/Z_10 , 
        \U3/U119/Z_9 , \U3/U119/Z_8 , n15364, n15365, n15366, n15367, 
        \U3/U105/Z_3 , \U3/U105/Z_2 , \U3/U105/Z_1 , \U3/U105/Z_0 }), .B({
        \U3/U118/Z_31 , \U3/U118/Z_30 , \U3/U118/Z_29 , \U3/U118/Z_28 , 
        \U3/U118/Z_27 , \U3/U118/Z_26 , \U3/U118/Z_25 , \U3/U118/Z_24 , 
        \U3/U118/Z_23 , \U3/U118/Z_22 , \U3/U118/Z_21 , \U3/U118/Z_20 , 
        \U3/U118/Z_19 , \U3/U118/Z_18 , \U3/U118/Z_17 , \U3/U118/Z_16 , 
        \U3/U118/Z_15 , \U3/U118/Z_14 , \U3/U118/Z_13 , \U3/U118/Z_12 , 
        \U3/U118/Z_11 , \U3/U118/Z_10 , \U3/U118/Z_9 , \U3/U118/Z_8 , n15371, 
        n15372, n15373, n15374, \U3/U106/Z_3 , n15375, \U3/U106/Z_1 , n15376}), 
        .LEQ(\U3/U107/Z_0 ), .TC(n15377), .LT_LE(N3336) );
  CannyEdge_DW01_addsub_16 r1044 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \U3/U81/Z_7 , \U3/U81/Z_6 , 
        \U3/U81/Z_5 , \U3/U81/Z_4 , \U3/U81/Z_3 , \U3/U81/Z_2 , \U3/U81/Z_1 , 
        \U3/U81/Z_0 }), .B({\U3/U82/Z_31 , \U3/U82/Z_30 , \U3/U82/Z_29 , 
        \U3/U82/Z_28 , \U3/U82/Z_27 , \U3/U82/Z_26 , \U3/U82/Z_25 , 
        \U3/U82/Z_24 , \U3/U82/Z_23 , \U3/U82/Z_22 , \U3/U82/Z_21 , 
        \U3/U82/Z_20 , \U3/U82/Z_19 , \U3/U82/Z_18 , \U3/U82/Z_17 , 
        \U3/U82/Z_16 , \U3/U82/Z_15 , \U3/U82/Z_14 , \U3/U82/Z_13 , 
        \U3/U82/Z_12 , \U3/U82/Z_11 , \U3/U82/Z_10 , \U3/U82/Z_9 , 
        \U3/U82/Z_8 , \U3/U82/Z_7 , \U3/U82/Z_6 , \U3/U82/Z_5 , \U3/U82/Z_4 , 
        \U3/U82/Z_3 , \U3/U82/Z_2 , \U3/U82/Z_1 , \U3/U82/Z_0 }), .CI(1'b0), 
        .ADD_SUB(n12467), .SUM({N2776, N2775, N2774, N2773, N2772, N2771, 
        N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, 
        N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, 
        N2750, N2749, N2748, N2747, N2746, N2648}) );
  CannyEdge_DW02_mult_24 r1023 ( .A({\U3/U64/Z_7 , \U3/U64/Z_6 , \U3/U64/Z_5 , 
        \U3/U64/Z_4 , \U3/U64/Z_3 , \U3/U64/Z_2 , \U3/U64/Z_1 , \U3/U64/Z_0 }), 
        .B({n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, n12477, 
        n12477, n12477, n12477, n12477, n12477, n12476, n12477, \U3/U65/Z_7 , 
        \U3/U65/Z_6 , \U3/U65/Z_5 , \U3/U65/Z_4 , \U3/U65/Z_3 , \U3/U65/Z_2 , 
        \U3/U65/Z_1 , \U3/U65/Z_0 }), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, N2267, N2266, 
        N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, 
        N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, 
        N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236})
         );
  OR2X2 U10044 ( .A(n12462), .B(n12570), .Y(n12461) );
  OR2X2 U10045 ( .A(IntSignal[1]), .B(IntSignal[0]), .Y(n12462) );
  AND2X2 U10046 ( .A(n13892), .B(n13893), .Y(n12463) );
  OR2X2 U10047 ( .A(n13058), .B(n14214), .Y(n12464) );
  OR2X2 U10048 ( .A(n13077), .B(n12537), .Y(n12465) );
  INVX2 U10049 ( .A(n12464), .Y(n12466) );
  INVX4 U10050 ( .A(n12463), .Y(n12467) );
  INVX4 U10051 ( .A(n12465), .Y(n12468) );
  INVX1 U10052 ( .A(n12554), .Y(n12469) );
  INVX4 U10053 ( .A(n12469), .Y(n12470) );
  INVX4 U10054 ( .A(n12462), .Y(n12471) );
  INVX1 U10055 ( .A(n12571), .Y(n12472) );
  INVX4 U10056 ( .A(n12472), .Y(n12473) );
  INVX4 U10057 ( .A(n15377), .Y(n14214) );
  INVX2 U10058 ( .A(n12905), .Y(n13034) );
  INVX2 U10059 ( .A(n13911), .Y(n13892) );
  BUFX2 U10060 ( .A(n13919), .Y(n12474) );
  INVX2 U10061 ( .A(n13905), .Y(n8303) );
  INVX2 U10062 ( .A(n13031), .Y(n12972) );
  AND2X2 U10063 ( .A(n12976), .B(IntSignal[1]), .Y(n12973) );
  AND2X2 U10064 ( .A(n13165), .B(n12473), .Y(n12976) );
  INVX2 U10065 ( .A(n12470), .Y(n15370) );
  BUFX4 U10066 ( .A(n15363), .Y(n12475) );
  INVX2 U10067 ( .A(n12475), .Y(n13893) );
  INVX4 U10068 ( .A(n12479), .Y(n12476) );
  INVX2 U10069 ( .A(n12478), .Y(n12477) );
  BUFX2 U10070 ( .A(n12461), .Y(n12483) );
  BUFX2 U10071 ( .A(n12461), .Y(n12485) );
  BUFX2 U10072 ( .A(n12461), .Y(n12484) );
  BUFX2 U10073 ( .A(n12461), .Y(n12478) );
  BUFX2 U10074 ( .A(n12461), .Y(n12479) );
  BUFX2 U10075 ( .A(n12461), .Y(n12488) );
  BUFX2 U10076 ( .A(n12461), .Y(n12487) );
  BUFX2 U10077 ( .A(n12489), .Y(n12480) );
  BUFX2 U10078 ( .A(n12461), .Y(n12481) );
  BUFX2 U10079 ( .A(n12489), .Y(n12482) );
  BUFX2 U10080 ( .A(n12461), .Y(n12486) );
  BUFX2 U10081 ( .A(n12461), .Y(n12489) );
  INVX1 U10082 ( .A(n12490), .Y(n15323) );
  MUX2X1 U10083 ( .B(InData[7]), .A(\regY[6][7] ), .S(n12491), .Y(n12490) );
  INVX1 U10084 ( .A(n12492), .Y(n15324) );
  MUX2X1 U10085 ( .B(InData[6]), .A(\regY[6][6] ), .S(n12491), .Y(n12492) );
  INVX1 U10086 ( .A(n12493), .Y(n15326) );
  AOI21X1 U10087 ( .A(n12494), .B(N976), .C(\U3/U100/Z_6 ), .Y(n12493) );
  INVX1 U10088 ( .A(n12495), .Y(n15329) );
  AOI22X1 U10089 ( .A(N2341), .B(n12476), .C(N2394), .D(n15370), .Y(n12495) );
  INVX1 U10090 ( .A(n12496), .Y(n15330) );
  AOI22X1 U10091 ( .A(N2340), .B(n12476), .C(N2393), .D(n15370), .Y(n12496) );
  INVX1 U10092 ( .A(n12497), .Y(n15331) );
  AOI22X1 U10093 ( .A(N2339), .B(n12476), .C(N2392), .D(n15370), .Y(n12497) );
  INVX1 U10094 ( .A(n12498), .Y(n15356) );
  AOI22X1 U10095 ( .A(N2338), .B(n12476), .C(N2391), .D(n15370), .Y(n12498) );
  INVX1 U10096 ( .A(n12499), .Y(n15357) );
  AOI22X1 U10097 ( .A(N2337), .B(n12476), .C(N2390), .D(n15370), .Y(n12499) );
  INVX1 U10098 ( .A(n12500), .Y(n15358) );
  AOI22X1 U10099 ( .A(N2336), .B(n12476), .C(N2389), .D(n15370), .Y(n12500) );
  INVX1 U10100 ( .A(n12501), .Y(n15359) );
  AOI22X1 U10101 ( .A(N2335), .B(n12476), .C(N2388), .D(n15370), .Y(n12501) );
  INVX1 U10102 ( .A(n12502), .Y(n15360) );
  AOI22X1 U10103 ( .A(N2334), .B(n12476), .C(N2387), .D(n15370), .Y(n12502) );
  INVX1 U10104 ( .A(n12503), .Y(n15361) );
  AOI22X1 U10105 ( .A(N2333), .B(n12476), .C(N2386), .D(n15370), .Y(n12503) );
  INVX1 U10106 ( .A(n12504), .Y(n15362) );
  AOI22X1 U10107 ( .A(N2332), .B(n12476), .C(N2385), .D(n15370), .Y(n12504) );
  INVX1 U10108 ( .A(n12505), .Y(n15364) );
  INVX1 U10109 ( .A(n12506), .Y(n15365) );
  INVX1 U10110 ( .A(n12507), .Y(n15366) );
  INVX1 U10111 ( .A(n12508), .Y(n15367) );
  OAI21X1 U10112 ( .A(n12509), .B(n12510), .C(n12511), .Y(n15368) );
  NAND3X1 U10113 ( .A(n12512), .B(n12513), .C(bCE), .Y(n12511) );
  INVX1 U10114 ( .A(n12514), .Y(n15371) );
  INVX1 U10115 ( .A(n12515), .Y(n15372) );
  INVX1 U10116 ( .A(n12516), .Y(n15373) );
  INVX1 U10117 ( .A(n12517), .Y(n15374) );
  INVX1 U10118 ( .A(N4438), .Y(n15464) );
  INVX1 U10119 ( .A(N4432), .Y(n15468) );
  INVX1 U10120 ( .A(N4468), .Y(n15846) );
  INVX1 U10121 ( .A(N4471), .Y(n15847) );
  INVX1 U10122 ( .A(N4474), .Y(n15848) );
  INVX1 U10123 ( .A(N4477), .Y(n15849) );
  INVX1 U10124 ( .A(N4480), .Y(n15850) );
  INVX1 U10125 ( .A(N4483), .Y(n15851) );
  INVX1 U10126 ( .A(N4486), .Y(n15852) );
  INVX1 U10127 ( .A(N4489), .Y(n15853) );
  MUX2X1 U10128 ( .B(n12518), .A(n12519), .S(n12520), .Y(n8322) );
  MUX2X1 U10129 ( .B(n12521), .A(n12522), .S(n12520), .Y(n8321) );
  MUX2X1 U10130 ( .B(n12523), .A(n12524), .S(n12520), .Y(n8320) );
  MUX2X1 U10131 ( .B(n12525), .A(n12526), .S(n12520), .Y(n8319) );
  MUX2X1 U10132 ( .B(n12527), .A(n12528), .S(n12520), .Y(n8318) );
  MUX2X1 U10133 ( .B(n12529), .A(n12530), .S(n12520), .Y(n8317) );
  MUX2X1 U10134 ( .B(n12531), .A(n12532), .S(n12520), .Y(n8316) );
  MUX2X1 U10135 ( .B(n12533), .A(n12534), .S(n12520), .Y(n8315) );
  NOR2X1 U10136 ( .A(n12535), .B(n12536), .Y(n12520) );
  INVX1 U10137 ( .A(n12537), .Y(n12536) );
  OAI21X1 U10138 ( .A(n12538), .B(n12539), .C(n12540), .Y(n8314) );
  INVX1 U10139 ( .A(n12541), .Y(n12540) );
  OAI22X1 U10140 ( .A(n12542), .B(n12543), .C(n12544), .D(n12545), .Y(n12541)
         );
  OR2X1 U10141 ( .A(n12546), .B(n12547), .Y(n12542) );
  INVX1 U10142 ( .A(n12548), .Y(n8291) );
  MUX2X1 U10143 ( .B(InData[1]), .A(\regY[6][1] ), .S(n12491), .Y(n12548) );
  INVX1 U10144 ( .A(n12549), .Y(n8289) );
  MUX2X1 U10145 ( .B(InData[3]), .A(\regY[6][3] ), .S(n12491), .Y(n12549) );
  INVX1 U10146 ( .A(n12550), .Y(n8288) );
  MUX2X1 U10147 ( .B(InData[4]), .A(\regY[6][4] ), .S(n12491), .Y(n12550) );
  INVX1 U10148 ( .A(n12551), .Y(n8287) );
  MUX2X1 U10149 ( .B(InData[5]), .A(\regY[6][5] ), .S(n12491), .Y(n12551) );
  OAI22X1 U10150 ( .A(n12552), .B(n12553), .C(n12470), .D(n12555), .Y(n5409)
         );
  OR2X1 U10151 ( .A(bCE), .B(dAddrRegRow[0]), .Y(n5398) );
  OR2X1 U10152 ( .A(bCE), .B(dAddrRegRow[1]), .Y(n5397) );
  AND2X1 U10153 ( .A(dAddrRegRow[2]), .B(n12556), .Y(n5396) );
  OAI21X1 U10154 ( .A(n15315), .B(n12557), .C(n12558), .Y(n5389) );
  INVX1 U10155 ( .A(N4469), .Y(n15315) );
  OAI21X1 U10156 ( .A(n15316), .B(n12557), .C(n12558), .Y(n5388) );
  INVX1 U10157 ( .A(N4472), .Y(n15316) );
  OAI21X1 U10158 ( .A(n15317), .B(n12557), .C(n12558), .Y(n5387) );
  INVX1 U10159 ( .A(N4475), .Y(n15317) );
  OAI21X1 U10160 ( .A(n15318), .B(n12557), .C(n12558), .Y(n5386) );
  INVX1 U10161 ( .A(N4478), .Y(n15318) );
  OAI21X1 U10162 ( .A(n15319), .B(n12557), .C(n12558), .Y(n5385) );
  INVX1 U10163 ( .A(N4481), .Y(n15319) );
  OAI21X1 U10164 ( .A(n15320), .B(n12557), .C(n12558), .Y(n5384) );
  INVX1 U10165 ( .A(N4484), .Y(n15320) );
  OAI21X1 U10166 ( .A(n15321), .B(n12557), .C(n12558), .Y(n5383) );
  INVX1 U10167 ( .A(N4487), .Y(n15321) );
  OAI21X1 U10168 ( .A(n15322), .B(n12557), .C(n12558), .Y(n5382) );
  NAND3X1 U10169 ( .A(n12559), .B(n12560), .C(n12557), .Y(n12558) );
  INVX1 U10170 ( .A(n12561), .Y(n12560) );
  NAND3X1 U10171 ( .A(n12562), .B(n12563), .C(n12564), .Y(n12559) );
  INVX1 U10172 ( .A(dReadReg[3]), .Y(n12563) );
  INVX1 U10173 ( .A(N4490), .Y(n15322) );
  OAI21X1 U10174 ( .A(n12509), .B(n12565), .C(n12566), .Y(n5381) );
  NAND3X1 U10175 ( .A(n12567), .B(n12513), .C(bCE), .Y(n12566) );
  OAI21X1 U10176 ( .A(OPMode[2]), .B(n12462), .C(n12568), .Y(n12567) );
  AND2X1 U10177 ( .A(bCE), .B(n12569), .Y(n12509) );
  OAI21X1 U10178 ( .A(n15377), .B(n12570), .C(n12513), .Y(n12569) );
  OAI21X1 U10179 ( .A(n15378), .B(n12473), .C(n12572), .Y(n5379) );
  INVX1 U10180 ( .A(N4466), .Y(n15378) );
  OAI21X1 U10181 ( .A(n15379), .B(n12473), .C(n12572), .Y(n5378) );
  INVX1 U10182 ( .A(N4463), .Y(n15379) );
  OAI21X1 U10183 ( .A(n15380), .B(n12473), .C(n12572), .Y(n5377) );
  INVX1 U10184 ( .A(N4460), .Y(n15380) );
  OAI21X1 U10185 ( .A(n15381), .B(n12473), .C(n12572), .Y(n5376) );
  INVX1 U10186 ( .A(N4457), .Y(n15381) );
  OAI21X1 U10187 ( .A(n15382), .B(n12473), .C(n12572), .Y(n5375) );
  INVX1 U10188 ( .A(N4454), .Y(n15382) );
  OAI21X1 U10189 ( .A(n15383), .B(n12473), .C(n12572), .Y(n5374) );
  INVX1 U10190 ( .A(N4451), .Y(n15383) );
  OAI21X1 U10191 ( .A(n15384), .B(n12473), .C(n12572), .Y(n5373) );
  INVX1 U10192 ( .A(N4448), .Y(n15384) );
  OAI21X1 U10193 ( .A(n15385), .B(n12473), .C(n12572), .Y(n5372) );
  INVX1 U10194 ( .A(N4445), .Y(n15385) );
  OAI21X1 U10195 ( .A(n15386), .B(n12473), .C(n12572), .Y(n5371) );
  INVX1 U10196 ( .A(N4373), .Y(n15386) );
  OAI21X1 U10197 ( .A(n15387), .B(n12473), .C(n12572), .Y(n5370) );
  INVX1 U10198 ( .A(N4376), .Y(n15387) );
  OAI21X1 U10199 ( .A(n15388), .B(n12473), .C(n12572), .Y(n5369) );
  INVX1 U10200 ( .A(N4379), .Y(n15388) );
  OAI21X1 U10201 ( .A(n15389), .B(n12473), .C(n12572), .Y(n5368) );
  INVX1 U10202 ( .A(N4382), .Y(n15389) );
  OAI21X1 U10203 ( .A(n15390), .B(n12473), .C(n12572), .Y(n5367) );
  INVX1 U10204 ( .A(N4385), .Y(n15390) );
  OAI21X1 U10205 ( .A(n15391), .B(n12473), .C(n12572), .Y(n5366) );
  INVX1 U10206 ( .A(N4388), .Y(n15391) );
  OAI21X1 U10207 ( .A(n15392), .B(n12473), .C(n12572), .Y(n5365) );
  INVX1 U10208 ( .A(N4391), .Y(n15392) );
  OAI21X1 U10209 ( .A(n15393), .B(n12473), .C(n12572), .Y(n5364) );
  NAND2X1 U10210 ( .A(n12473), .B(n12573), .Y(n12572) );
  INVX1 U10211 ( .A(N4394), .Y(n15393) );
  AOI21X1 U10212 ( .A(n15394), .B(n12574), .C(n12575), .Y(n5363) );
  INVX1 U10213 ( .A(N4502), .Y(n15394) );
  MUX2X1 U10214 ( .B(n12576), .A(n12577), .S(n12578), .Y(n5362) );
  MUX2X1 U10215 ( .B(n12579), .A(n12580), .S(n12578), .Y(n5361) );
  MUX2X1 U10216 ( .B(n12581), .A(n12582), .S(n12578), .Y(n5360) );
  MUX2X1 U10217 ( .B(n12583), .A(n12584), .S(n12578), .Y(n5359) );
  MUX2X1 U10218 ( .B(n12585), .A(n12586), .S(n12578), .Y(n5358) );
  MUX2X1 U10219 ( .B(n12587), .A(n12588), .S(n12578), .Y(n5357) );
  MUX2X1 U10220 ( .B(n12589), .A(n12590), .S(n12578), .Y(n5356) );
  MUX2X1 U10221 ( .B(n12591), .A(n12592), .S(n12578), .Y(n5355) );
  OAI22X1 U10222 ( .A(n12593), .B(n12594), .C(n12595), .D(n12596), .Y(n12578)
         );
  MUX2X1 U10223 ( .B(n12582), .A(n12597), .S(n12598), .Y(n5354) );
  MUX2X1 U10224 ( .B(n12584), .A(n12599), .S(n12598), .Y(n5353) );
  MUX2X1 U10225 ( .B(n12586), .A(n12600), .S(n12598), .Y(n5352) );
  MUX2X1 U10226 ( .B(n12588), .A(n12601), .S(n12598), .Y(n5351) );
  MUX2X1 U10227 ( .B(n12590), .A(n12602), .S(n12598), .Y(n5350) );
  MUX2X1 U10228 ( .B(n12592), .A(n12603), .S(n12598), .Y(n5349) );
  MUX2X1 U10229 ( .B(n12580), .A(n12604), .S(n12598), .Y(n5348) );
  MUX2X1 U10230 ( .B(n12577), .A(n12605), .S(n12598), .Y(n5347) );
  AOI22X1 U10231 ( .A(n12606), .B(n12607), .C(n12608), .D(n12609), .Y(n12598)
         );
  MUX2X1 U10232 ( .B(n12610), .A(n12592), .S(n12611), .Y(n5346) );
  MUX2X1 U10233 ( .B(n12612), .A(n12590), .S(n12611), .Y(n5345) );
  MUX2X1 U10234 ( .B(n12613), .A(n12588), .S(n12611), .Y(n5344) );
  MUX2X1 U10235 ( .B(n12614), .A(n12586), .S(n12611), .Y(n5343) );
  MUX2X1 U10236 ( .B(n12615), .A(n12584), .S(n12611), .Y(n5342) );
  MUX2X1 U10237 ( .B(n12616), .A(n12582), .S(n12611), .Y(n5341) );
  MUX2X1 U10238 ( .B(n12617), .A(n12580), .S(n12611), .Y(n5340) );
  MUX2X1 U10239 ( .B(n12618), .A(n12577), .S(n12611), .Y(n5339) );
  OAI22X1 U10240 ( .A(n12593), .B(n12619), .C(n12595), .D(n12620), .Y(n12611)
         );
  MUX2X1 U10241 ( .B(n15395), .A(n12621), .S(n12622), .Y(n5338) );
  INVX1 U10242 ( .A(N4081), .Y(n15395) );
  OAI21X1 U10243 ( .A(n15396), .B(n12622), .C(n12623), .Y(n5337) );
  INVX1 U10244 ( .A(N4082), .Y(n15396) );
  OAI21X1 U10245 ( .A(n15397), .B(n12622), .C(n12623), .Y(n5336) );
  INVX1 U10246 ( .A(N4061), .Y(n15397) );
  MUX2X1 U10247 ( .B(n15398), .A(n12624), .S(n12622), .Y(n5335) );
  INVX1 U10248 ( .A(N4060), .Y(n15398) );
  OAI21X1 U10249 ( .A(n15399), .B(n12622), .C(n12623), .Y(n5334) );
  INVX1 U10250 ( .A(N4064), .Y(n15399) );
  MUX2X1 U10251 ( .B(n15400), .A(n12625), .S(n12622), .Y(n5333) );
  INVX1 U10252 ( .A(N4063), .Y(n15400) );
  OAI21X1 U10253 ( .A(n15401), .B(n12622), .C(n12623), .Y(n5332) );
  INVX1 U10254 ( .A(N4067), .Y(n15401) );
  MUX2X1 U10255 ( .B(n15402), .A(n12626), .S(n12622), .Y(n5331) );
  INVX1 U10256 ( .A(N4066), .Y(n15402) );
  OAI21X1 U10257 ( .A(n15403), .B(n12622), .C(n12623), .Y(n5330) );
  INVX1 U10258 ( .A(N4070), .Y(n15403) );
  MUX2X1 U10259 ( .B(n15404), .A(n12627), .S(n12622), .Y(n5329) );
  INVX1 U10260 ( .A(N4069), .Y(n15404) );
  OAI21X1 U10261 ( .A(n15405), .B(n12622), .C(n12623), .Y(n5328) );
  INVX1 U10262 ( .A(N4073), .Y(n15405) );
  MUX2X1 U10263 ( .B(n15406), .A(n12628), .S(n12622), .Y(n5327) );
  INVX1 U10264 ( .A(N4072), .Y(n15406) );
  OAI21X1 U10265 ( .A(n15407), .B(n12622), .C(n12623), .Y(n5326) );
  INVX1 U10266 ( .A(N4076), .Y(n15407) );
  MUX2X1 U10267 ( .B(n15408), .A(n12629), .S(n12622), .Y(n5325) );
  INVX1 U10268 ( .A(N4075), .Y(n15408) );
  OAI21X1 U10269 ( .A(n15409), .B(n12622), .C(n12623), .Y(n5324) );
  NAND2X1 U10270 ( .A(n12630), .B(n12622), .Y(n12623) );
  INVX1 U10271 ( .A(N4079), .Y(n15409) );
  MUX2X1 U10272 ( .B(n15410), .A(n12631), .S(n12622), .Y(n5323) );
  AND2X1 U10273 ( .A(n12632), .B(n12633), .Y(n12622) );
  INVX1 U10274 ( .A(N4078), .Y(n15410) );
  MUX2X1 U10275 ( .B(n15411), .A(n12621), .S(n12634), .Y(n5322) );
  INVX1 U10276 ( .A(N3793), .Y(n15411) );
  OAI21X1 U10277 ( .A(n15412), .B(n12634), .C(n12635), .Y(n5321) );
  INVX1 U10278 ( .A(N3794), .Y(n15412) );
  MUX2X1 U10279 ( .B(n15413), .A(n12631), .S(n12634), .Y(n5320) );
  INVX1 U10280 ( .A(N3790), .Y(n15413) );
  OAI21X1 U10281 ( .A(n15414), .B(n12634), .C(n12635), .Y(n5319) );
  INVX1 U10282 ( .A(N3791), .Y(n15414) );
  MUX2X1 U10283 ( .B(n15415), .A(n12629), .S(n12634), .Y(n5318) );
  INVX1 U10284 ( .A(N3787), .Y(n15415) );
  OAI21X1 U10285 ( .A(n15416), .B(n12634), .C(n12635), .Y(n5317) );
  INVX1 U10286 ( .A(N3788), .Y(n15416) );
  MUX2X1 U10287 ( .B(n15417), .A(n12628), .S(n12634), .Y(n5316) );
  INVX1 U10288 ( .A(N3784), .Y(n15417) );
  OAI21X1 U10289 ( .A(n15418), .B(n12634), .C(n12635), .Y(n5315) );
  INVX1 U10290 ( .A(N3785), .Y(n15418) );
  OAI21X1 U10291 ( .A(n15419), .B(n12634), .C(n12635), .Y(n5314) );
  INVX1 U10292 ( .A(N3773), .Y(n15419) );
  MUX2X1 U10293 ( .B(n15420), .A(n12624), .S(n12634), .Y(n5313) );
  INVX1 U10294 ( .A(N3772), .Y(n15420) );
  OAI21X1 U10295 ( .A(n15421), .B(n12634), .C(n12635), .Y(n5312) );
  INVX1 U10296 ( .A(N3776), .Y(n15421) );
  MUX2X1 U10297 ( .B(n15422), .A(n12625), .S(n12634), .Y(n5311) );
  INVX1 U10298 ( .A(N3775), .Y(n15422) );
  OAI21X1 U10299 ( .A(n15423), .B(n12634), .C(n12635), .Y(n5310) );
  INVX1 U10300 ( .A(N3779), .Y(n15423) );
  MUX2X1 U10301 ( .B(n15424), .A(n12626), .S(n12634), .Y(n5309) );
  INVX1 U10302 ( .A(N3778), .Y(n15424) );
  OAI21X1 U10303 ( .A(n15425), .B(n12634), .C(n12635), .Y(n5308) );
  NAND2X1 U10304 ( .A(n12634), .B(n12630), .Y(n12635) );
  INVX1 U10305 ( .A(N3782), .Y(n15425) );
  MUX2X1 U10306 ( .B(n15426), .A(n12627), .S(n12634), .Y(n5307) );
  AND2X1 U10307 ( .A(n12636), .B(n12607), .Y(n12634) );
  INVX1 U10308 ( .A(N3781), .Y(n15426) );
  OAI21X1 U10309 ( .A(n12538), .B(n12637), .C(n12638), .Y(n5297) );
  INVX1 U10310 ( .A(dy[1]), .Y(n12637) );
  OR2X1 U10311 ( .A(n12639), .B(n12640), .Y(n5296) );
  OAI22X1 U10312 ( .A(n15427), .B(n12538), .C(n12544), .D(n12641), .Y(n12640)
         );
  INVX1 U10313 ( .A(N4501), .Y(n15427) );
  OAI21X1 U10314 ( .A(n12547), .B(n12642), .C(n12638), .Y(n12639) );
  OR2X1 U10315 ( .A(n12643), .B(n12644), .Y(n5295) );
  OAI22X1 U10316 ( .A(n15428), .B(n12538), .C(n12544), .D(n12642), .Y(n12644)
         );
  NAND2X1 U10317 ( .A(n12538), .B(OPMode[0]), .Y(n12544) );
  INVX1 U10318 ( .A(N4495), .Y(n15428) );
  OAI21X1 U10319 ( .A(n12547), .B(n12641), .C(n12638), .Y(n12643) );
  NAND2X1 U10320 ( .A(n12538), .B(n12645), .Y(n12638) );
  NAND2X1 U10321 ( .A(n12538), .B(n12646), .Y(n12547) );
  AOI21X1 U10322 ( .A(n15429), .B(n12574), .C(n12575), .Y(n5294) );
  INVX1 U10323 ( .A(n12647), .Y(n12575) );
  OAI21X1 U10324 ( .A(n12645), .B(n12648), .C(n12538), .Y(n12647) );
  INVX1 U10325 ( .A(n12574), .Y(n12538) );
  NAND2X1 U10326 ( .A(n12642), .B(n12641), .Y(n12648) );
  OR2X1 U10327 ( .A(n12649), .B(n12650), .Y(n12641) );
  NAND3X1 U10328 ( .A(\regY[6][4] ), .B(\regY[6][3] ), .C(n12651), .Y(n12650)
         );
  NAND3X1 U10329 ( .A(\regY[6][6] ), .B(n12652), .C(\regY[6][1] ), .Y(n12649)
         );
  INVX1 U10330 ( .A(\regY[6][5] ), .Y(n12652) );
  NAND3X1 U10331 ( .A(n12653), .B(n12654), .C(n12651), .Y(n12642) );
  INVX1 U10332 ( .A(n12655), .Y(n12651) );
  NAND3X1 U10333 ( .A(n12656), .B(n12657), .C(n12658), .Y(n12655) );
  INVX1 U10334 ( .A(n12546), .Y(n12653) );
  OAI21X1 U10335 ( .A(n12546), .B(n12543), .C(n12545), .Y(n12645) );
  OR2X1 U10336 ( .A(n12659), .B(n12660), .Y(n12545) );
  NAND3X1 U10337 ( .A(\regY[6][5] ), .B(\regY[6][3] ), .C(n12661), .Y(n12660)
         );
  NOR2X1 U10338 ( .A(n12658), .B(n12656), .Y(n12661) );
  INVX1 U10339 ( .A(\regY[6][2] ), .Y(n12656) );
  NAND3X1 U10340 ( .A(n12654), .B(n12662), .C(n12663), .Y(n12659) );
  NOR2X1 U10341 ( .A(\regY[6][7] ), .B(\regY[6][6] ), .Y(n12663) );
  INVX1 U10342 ( .A(\regY[6][1] ), .Y(n12654) );
  NAND3X1 U10343 ( .A(\regY[6][2] ), .B(\regY[6][1] ), .C(n12664), .Y(n12543)
         );
  NOR2X1 U10344 ( .A(n12657), .B(n12658), .Y(n12664) );
  INVX1 U10345 ( .A(\regY[6][0] ), .Y(n12658) );
  INVX1 U10346 ( .A(\regY[6][7] ), .Y(n12657) );
  NAND3X1 U10347 ( .A(n12665), .B(n12662), .C(n12666), .Y(n12546) );
  NOR2X1 U10348 ( .A(\regY[6][6] ), .B(\regY[6][5] ), .Y(n12666) );
  INVX1 U10349 ( .A(\regY[6][4] ), .Y(n12662) );
  INVX1 U10350 ( .A(\regY[6][3] ), .Y(n12665) );
  NAND3X1 U10351 ( .A(n12471), .B(n12667), .C(n12668), .Y(n12574) );
  INVX1 U10352 ( .A(N4496), .Y(n15429) );
  MUX2X1 U10353 ( .B(n12669), .A(n12577), .S(n12670), .Y(n5293) );
  MUX2X1 U10354 ( .B(n12671), .A(n12580), .S(n12670), .Y(n5292) );
  MUX2X1 U10355 ( .B(n12672), .A(n12582), .S(n12670), .Y(n5291) );
  MUX2X1 U10356 ( .B(n12673), .A(n12584), .S(n12670), .Y(n5290) );
  MUX2X1 U10357 ( .B(n12674), .A(n12586), .S(n12670), .Y(n5289) );
  MUX2X1 U10358 ( .B(n12675), .A(n12588), .S(n12670), .Y(n5288) );
  MUX2X1 U10359 ( .B(n12676), .A(n12590), .S(n12670), .Y(n5287) );
  MUX2X1 U10360 ( .B(n12677), .A(n12592), .S(n12670), .Y(n5286) );
  OAI22X1 U10361 ( .A(n12678), .B(n12679), .C(n12680), .D(n12681), .Y(n12670)
         );
  OAI21X1 U10362 ( .A(n12682), .B(n12683), .C(n15369), .Y(n12681) );
  OAI21X1 U10363 ( .A(n12678), .B(n12684), .C(N2777), .Y(n12683) );
  OAI21X1 U10364 ( .A(n12685), .B(n12686), .C(n12687), .Y(n12682) );
  NAND2X1 U10365 ( .A(n12688), .B(n12689), .Y(n12686) );
  MUX2X1 U10366 ( .B(n12577), .A(n12690), .S(n12691), .Y(n5285) );
  MUX2X1 U10367 ( .B(n12580), .A(n12692), .S(n12691), .Y(n5284) );
  MUX2X1 U10368 ( .B(n12582), .A(n12693), .S(n12691), .Y(n5283) );
  MUX2X1 U10369 ( .B(n12584), .A(n12694), .S(n12691), .Y(n5282) );
  MUX2X1 U10370 ( .B(n12586), .A(n12695), .S(n12691), .Y(n5281) );
  MUX2X1 U10371 ( .B(n12588), .A(n12696), .S(n12691), .Y(n5280) );
  MUX2X1 U10372 ( .B(n12590), .A(n12697), .S(n12691), .Y(n5279) );
  MUX2X1 U10373 ( .B(n12592), .A(n12698), .S(n12691), .Y(n5278) );
  AOI22X1 U10374 ( .A(n12606), .B(n12699), .C(n12608), .D(n12700), .Y(n12691)
         );
  MUX2X1 U10375 ( .B(n12577), .A(n12701), .S(n12702), .Y(n5277) );
  MUX2X1 U10376 ( .B(n12580), .A(n12703), .S(n12702), .Y(n5276) );
  MUX2X1 U10377 ( .B(n12582), .A(n12704), .S(n12702), .Y(n5275) );
  MUX2X1 U10378 ( .B(n12584), .A(n12705), .S(n12702), .Y(n5274) );
  MUX2X1 U10379 ( .B(n12586), .A(n12706), .S(n12702), .Y(n5273) );
  MUX2X1 U10380 ( .B(n12588), .A(n12707), .S(n12702), .Y(n5272) );
  MUX2X1 U10381 ( .B(n12590), .A(n12708), .S(n12702), .Y(n5271) );
  MUX2X1 U10382 ( .B(n12592), .A(n12709), .S(n12702), .Y(n5270) );
  AOI22X1 U10383 ( .A(n12606), .B(n12710), .C(n12608), .D(n12711), .Y(n12702)
         );
  MUX2X1 U10384 ( .B(n12577), .A(n12712), .S(n12713), .Y(n5269) );
  MUX2X1 U10385 ( .B(n12580), .A(n12714), .S(n12713), .Y(n5268) );
  MUX2X1 U10386 ( .B(n12582), .A(n12715), .S(n12713), .Y(n5267) );
  MUX2X1 U10387 ( .B(n12584), .A(n12716), .S(n12713), .Y(n5266) );
  MUX2X1 U10388 ( .B(n12586), .A(n12717), .S(n12713), .Y(n5265) );
  MUX2X1 U10389 ( .B(n12588), .A(n12718), .S(n12713), .Y(n5264) );
  MUX2X1 U10390 ( .B(n12590), .A(n12719), .S(n12713), .Y(n5263) );
  MUX2X1 U10391 ( .B(n12592), .A(n12720), .S(n12713), .Y(n5262) );
  AOI22X1 U10392 ( .A(n12606), .B(n12721), .C(n12608), .D(n12722), .Y(n12713)
         );
  INVX1 U10393 ( .A(n12723), .Y(n12721) );
  MUX2X1 U10394 ( .B(n12577), .A(n12724), .S(n12725), .Y(n5261) );
  MUX2X1 U10395 ( .B(n12580), .A(n12726), .S(n12725), .Y(n5260) );
  MUX2X1 U10396 ( .B(n12582), .A(n12727), .S(n12725), .Y(n5259) );
  MUX2X1 U10397 ( .B(n12584), .A(n12728), .S(n12725), .Y(n5258) );
  MUX2X1 U10398 ( .B(n12586), .A(n12729), .S(n12725), .Y(n5257) );
  MUX2X1 U10399 ( .B(n12588), .A(n12730), .S(n12725), .Y(n5256) );
  MUX2X1 U10400 ( .B(n12590), .A(n12731), .S(n12725), .Y(n5255) );
  MUX2X1 U10401 ( .B(n12592), .A(n12732), .S(n12725), .Y(n5254) );
  AOI22X1 U10402 ( .A(n12606), .B(n12733), .C(n12608), .D(n12734), .Y(n12725)
         );
  INVX1 U10403 ( .A(n12735), .Y(n12733) );
  MUX2X1 U10404 ( .B(n12577), .A(n12736), .S(n12737), .Y(n5253) );
  MUX2X1 U10405 ( .B(n12580), .A(n12738), .S(n12737), .Y(n5252) );
  MUX2X1 U10406 ( .B(n12582), .A(n12739), .S(n12737), .Y(n5251) );
  MUX2X1 U10407 ( .B(n12584), .A(n12740), .S(n12737), .Y(n5250) );
  MUX2X1 U10408 ( .B(n12586), .A(n12741), .S(n12737), .Y(n5249) );
  MUX2X1 U10409 ( .B(n12588), .A(n12742), .S(n12737), .Y(n5248) );
  MUX2X1 U10410 ( .B(n12590), .A(n12743), .S(n12737), .Y(n5247) );
  MUX2X1 U10411 ( .B(n12592), .A(n12744), .S(n12737), .Y(n5246) );
  AOI22X1 U10412 ( .A(n12606), .B(n12745), .C(n12608), .D(n12746), .Y(n12737)
         );
  MUX2X1 U10413 ( .B(n12577), .A(n12747), .S(n12748), .Y(n5245) );
  MUX2X1 U10414 ( .B(n12580), .A(n12749), .S(n12748), .Y(n5244) );
  MUX2X1 U10415 ( .B(n12582), .A(n12750), .S(n12748), .Y(n5243) );
  MUX2X1 U10416 ( .B(n12584), .A(n12751), .S(n12748), .Y(n5242) );
  MUX2X1 U10417 ( .B(n12586), .A(n12752), .S(n12748), .Y(n5241) );
  MUX2X1 U10418 ( .B(n12588), .A(n12753), .S(n12748), .Y(n5240) );
  MUX2X1 U10419 ( .B(n12590), .A(n12754), .S(n12748), .Y(n5239) );
  MUX2X1 U10420 ( .B(n12592), .A(n12755), .S(n12748), .Y(n5238) );
  AOI22X1 U10421 ( .A(n12606), .B(n12756), .C(n12757), .D(n12608), .Y(n12748)
         );
  NOR2X1 U10422 ( .A(n12758), .B(n12759), .Y(n12608) );
  MUX2X1 U10423 ( .B(n12577), .A(n12760), .S(n12761), .Y(n5237) );
  MUX2X1 U10424 ( .B(n12580), .A(n12762), .S(n12761), .Y(n5236) );
  MUX2X1 U10425 ( .B(n12582), .A(n12763), .S(n12761), .Y(n5235) );
  MUX2X1 U10426 ( .B(n12584), .A(n12764), .S(n12761), .Y(n5234) );
  MUX2X1 U10427 ( .B(n12586), .A(n12765), .S(n12761), .Y(n5233) );
  MUX2X1 U10428 ( .B(n12588), .A(n12766), .S(n12761), .Y(n5232) );
  MUX2X1 U10429 ( .B(n12590), .A(n12767), .S(n12761), .Y(n5231) );
  MUX2X1 U10430 ( .B(n12592), .A(n12768), .S(n12761), .Y(n5230) );
  AOI22X1 U10431 ( .A(n12606), .B(n12769), .C(n12770), .D(n12609), .Y(n12761)
         );
  MUX2X1 U10432 ( .B(n12577), .A(n12771), .S(n12772), .Y(n5229) );
  MUX2X1 U10433 ( .B(n12580), .A(n12773), .S(n12772), .Y(n5228) );
  MUX2X1 U10434 ( .B(n12582), .A(n12774), .S(n12772), .Y(n5227) );
  MUX2X1 U10435 ( .B(n12584), .A(n12775), .S(n12772), .Y(n5226) );
  MUX2X1 U10436 ( .B(n12586), .A(n12776), .S(n12772), .Y(n5225) );
  MUX2X1 U10437 ( .B(n12588), .A(n12777), .S(n12772), .Y(n5224) );
  MUX2X1 U10438 ( .B(n12590), .A(n12778), .S(n12772), .Y(n5223) );
  MUX2X1 U10439 ( .B(n12592), .A(n12779), .S(n12772), .Y(n5222) );
  AOI22X1 U10440 ( .A(n12780), .B(n12781), .C(n12770), .D(n12700), .Y(n12772)
         );
  MUX2X1 U10441 ( .B(n12577), .A(n12782), .S(n12783), .Y(n5221) );
  MUX2X1 U10442 ( .B(n12580), .A(n12784), .S(n12783), .Y(n5220) );
  MUX2X1 U10443 ( .B(n12582), .A(n12785), .S(n12783), .Y(n5219) );
  MUX2X1 U10444 ( .B(n12584), .A(n12786), .S(n12783), .Y(n5218) );
  MUX2X1 U10445 ( .B(n12586), .A(n12787), .S(n12783), .Y(n5217) );
  INVX1 U10446 ( .A(\regX[16][4] ), .Y(n12787) );
  MUX2X1 U10447 ( .B(n12588), .A(n12788), .S(n12783), .Y(n5216) );
  INVX1 U10448 ( .A(\regX[16][5] ), .Y(n12788) );
  MUX2X1 U10449 ( .B(n12590), .A(n12789), .S(n12783), .Y(n5215) );
  INVX1 U10450 ( .A(\regX[16][6] ), .Y(n12789) );
  MUX2X1 U10451 ( .B(n12592), .A(n12790), .S(n12783), .Y(n5214) );
  AOI22X1 U10452 ( .A(n12606), .B(n12791), .C(n12609), .D(n12792), .Y(n12783)
         );
  INVX1 U10453 ( .A(\regX[16][7] ), .Y(n12790) );
  MUX2X1 U10454 ( .B(n12577), .A(n12793), .S(n12794), .Y(n5213) );
  MUX2X1 U10455 ( .B(n12580), .A(n12795), .S(n12794), .Y(n5212) );
  MUX2X1 U10456 ( .B(n12582), .A(n12796), .S(n12794), .Y(n5211) );
  MUX2X1 U10457 ( .B(n12584), .A(n12797), .S(n12794), .Y(n5210) );
  MUX2X1 U10458 ( .B(n12586), .A(n12798), .S(n12794), .Y(n5209) );
  MUX2X1 U10459 ( .B(n12588), .A(n12799), .S(n12794), .Y(n5208) );
  MUX2X1 U10460 ( .B(n12590), .A(n12800), .S(n12794), .Y(n5207) );
  MUX2X1 U10461 ( .B(n12592), .A(n12801), .S(n12794), .Y(n5206) );
  AOI22X1 U10462 ( .A(n12802), .B(n12803), .C(n12700), .D(n12792), .Y(n12794)
         );
  MUX2X1 U10463 ( .B(n12804), .A(n12577), .S(n12805), .Y(n5205) );
  MUX2X1 U10464 ( .B(n12806), .A(n12580), .S(n12805), .Y(n5204) );
  MUX2X1 U10465 ( .B(n12807), .A(n12582), .S(n12805), .Y(n5203) );
  MUX2X1 U10466 ( .B(n12808), .A(n12584), .S(n12805), .Y(n5202) );
  MUX2X1 U10467 ( .B(n12809), .A(n12586), .S(n12805), .Y(n5201) );
  MUX2X1 U10468 ( .B(n12810), .A(n12588), .S(n12805), .Y(n5200) );
  MUX2X1 U10469 ( .B(n12811), .A(n12590), .S(n12805), .Y(n5199) );
  MUX2X1 U10470 ( .B(n12812), .A(n12592), .S(n12805), .Y(n5198) );
  OAI21X1 U10471 ( .A(n12813), .B(n12814), .C(n12815), .Y(n12805) );
  NAND3X1 U10472 ( .A(n12816), .B(n12606), .C(n12817), .Y(n12815) );
  NAND2X1 U10473 ( .A(n12609), .B(n12818), .Y(n12814) );
  NAND2X1 U10474 ( .A(n12819), .B(n12820), .Y(n12813) );
  MUX2X1 U10475 ( .B(n12577), .A(n12821), .S(n12822), .Y(n5197) );
  MUX2X1 U10476 ( .B(n12580), .A(n12823), .S(n12822), .Y(n5196) );
  MUX2X1 U10477 ( .B(n12582), .A(n12824), .S(n12822), .Y(n5195) );
  MUX2X1 U10478 ( .B(n12584), .A(n12825), .S(n12822), .Y(n5194) );
  MUX2X1 U10479 ( .B(n12586), .A(n12826), .S(n12822), .Y(n5193) );
  MUX2X1 U10480 ( .B(n12588), .A(n12827), .S(n12822), .Y(n5192) );
  MUX2X1 U10481 ( .B(n12590), .A(n12828), .S(n12822), .Y(n5191) );
  MUX2X1 U10482 ( .B(n12592), .A(n12829), .S(n12822), .Y(n5190) );
  AOI22X1 U10483 ( .A(n12780), .B(n12830), .C(n12770), .D(n12831), .Y(n12822)
         );
  MUX2X1 U10484 ( .B(n12577), .A(n12832), .S(n12833), .Y(n5189) );
  MUX2X1 U10485 ( .B(n12580), .A(n12834), .S(n12833), .Y(n5188) );
  MUX2X1 U10486 ( .B(n12582), .A(n12835), .S(n12833), .Y(n5187) );
  MUX2X1 U10487 ( .B(n12584), .A(n12836), .S(n12833), .Y(n5186) );
  MUX2X1 U10488 ( .B(n12586), .A(n12837), .S(n12833), .Y(n5185) );
  MUX2X1 U10489 ( .B(n12588), .A(n12838), .S(n12833), .Y(n5184) );
  MUX2X1 U10490 ( .B(n12590), .A(n12839), .S(n12833), .Y(n5183) );
  MUX2X1 U10491 ( .B(n12592), .A(n12840), .S(n12833), .Y(n5182) );
  AOI22X1 U10492 ( .A(n12802), .B(n12841), .C(n12831), .D(n12792), .Y(n12833)
         );
  MUX2X1 U10493 ( .B(n12577), .A(n12842), .S(n12843), .Y(n5181) );
  MUX2X1 U10494 ( .B(n12580), .A(n12844), .S(n12843), .Y(n5180) );
  MUX2X1 U10495 ( .B(n12582), .A(n12845), .S(n12843), .Y(n5179) );
  MUX2X1 U10496 ( .B(n12584), .A(n12846), .S(n12843), .Y(n5178) );
  MUX2X1 U10497 ( .B(n12586), .A(n12847), .S(n12843), .Y(n5177) );
  MUX2X1 U10498 ( .B(n12588), .A(n12848), .S(n12843), .Y(n5176) );
  MUX2X1 U10499 ( .B(n12590), .A(n12849), .S(n12843), .Y(n5175) );
  MUX2X1 U10500 ( .B(n12592), .A(n12850), .S(n12843), .Y(n5174) );
  AOI22X1 U10501 ( .A(n12802), .B(n12851), .C(n12757), .D(n12792), .Y(n12843)
         );
  MUX2X1 U10502 ( .B(n12577), .A(n12852), .S(n12853), .Y(n5173) );
  MUX2X1 U10503 ( .B(n12580), .A(n12854), .S(n12853), .Y(n5172) );
  MUX2X1 U10504 ( .B(n12582), .A(n12855), .S(n12853), .Y(n5171) );
  MUX2X1 U10505 ( .B(n12584), .A(n12856), .S(n12853), .Y(n5170) );
  MUX2X1 U10506 ( .B(n12586), .A(n12857), .S(n12853), .Y(n5169) );
  MUX2X1 U10507 ( .B(n12588), .A(n12858), .S(n12853), .Y(n5168) );
  MUX2X1 U10508 ( .B(n12590), .A(n12859), .S(n12853), .Y(n5167) );
  MUX2X1 U10509 ( .B(n12592), .A(n12860), .S(n12853), .Y(n5166) );
  AOI22X1 U10510 ( .A(n12780), .B(n12632), .C(n12770), .D(n12734), .Y(n12853)
         );
  MUX2X1 U10511 ( .B(n12577), .A(n12861), .S(n12862), .Y(n5165) );
  MUX2X1 U10512 ( .B(n12580), .A(n12863), .S(n12862), .Y(n5164) );
  MUX2X1 U10513 ( .B(n12582), .A(n12864), .S(n12862), .Y(n5163) );
  MUX2X1 U10514 ( .B(n12584), .A(n12865), .S(n12862), .Y(n5162) );
  MUX2X1 U10515 ( .B(n12586), .A(n12866), .S(n12862), .Y(n5161) );
  MUX2X1 U10516 ( .B(n12588), .A(n12867), .S(n12862), .Y(n5160) );
  MUX2X1 U10517 ( .B(n12590), .A(n12868), .S(n12862), .Y(n5159) );
  MUX2X1 U10518 ( .B(n12592), .A(n12869), .S(n12862), .Y(n5158) );
  AOI22X1 U10519 ( .A(n12802), .B(n12870), .C(n12734), .D(n12792), .Y(n12862)
         );
  MUX2X1 U10520 ( .B(n12577), .A(n12871), .S(n12872), .Y(n5157) );
  MUX2X1 U10521 ( .B(n12580), .A(n12873), .S(n12872), .Y(n5156) );
  MUX2X1 U10522 ( .B(n12582), .A(n12874), .S(n12872), .Y(n5155) );
  MUX2X1 U10523 ( .B(n12584), .A(n12875), .S(n12872), .Y(n5154) );
  MUX2X1 U10524 ( .B(n12586), .A(n12876), .S(n12872), .Y(n5153) );
  MUX2X1 U10525 ( .B(n12588), .A(n12877), .S(n12872), .Y(n5152) );
  MUX2X1 U10526 ( .B(n12590), .A(n12878), .S(n12872), .Y(n5151) );
  MUX2X1 U10527 ( .B(n12592), .A(n12879), .S(n12872), .Y(n5150) );
  AOI22X1 U10528 ( .A(n12802), .B(n12880), .C(n12746), .D(n12792), .Y(n12872)
         );
  MUX2X1 U10529 ( .B(n12577), .A(n12881), .S(n12882), .Y(n5149) );
  MUX2X1 U10530 ( .B(n12580), .A(n12883), .S(n12882), .Y(n5148) );
  MUX2X1 U10531 ( .B(n12582), .A(n12884), .S(n12882), .Y(n5147) );
  MUX2X1 U10532 ( .B(n12584), .A(n12885), .S(n12882), .Y(n5146) );
  MUX2X1 U10533 ( .B(n12586), .A(n12886), .S(n12882), .Y(n5145) );
  MUX2X1 U10534 ( .B(n12588), .A(n12887), .S(n12882), .Y(n5144) );
  MUX2X1 U10535 ( .B(n12590), .A(n12888), .S(n12882), .Y(n5143) );
  MUX2X1 U10536 ( .B(n12592), .A(n12889), .S(n12882), .Y(n5142) );
  AOI22X1 U10537 ( .A(n12780), .B(n12890), .C(n12770), .D(n12711), .Y(n12882)
         );
  MUX2X1 U10538 ( .B(n12577), .A(n12891), .S(n12892), .Y(n5141) );
  MUX2X1 U10539 ( .B(n12580), .A(n12893), .S(n12892), .Y(n5140) );
  MUX2X1 U10540 ( .B(n12582), .A(n12894), .S(n12892), .Y(n5139) );
  MUX2X1 U10541 ( .B(n12584), .A(n12895), .S(n12892), .Y(n5138) );
  MUX2X1 U10542 ( .B(n12586), .A(n12896), .S(n12892), .Y(n5137) );
  MUX2X1 U10543 ( .B(n12588), .A(n12897), .S(n12892), .Y(n5136) );
  MUX2X1 U10544 ( .B(n12590), .A(n12898), .S(n12892), .Y(n5135) );
  MUX2X1 U10545 ( .B(n12592), .A(n12899), .S(n12892), .Y(n5134) );
  AOI22X1 U10546 ( .A(n12780), .B(n12900), .C(n12770), .D(n12722), .Y(n12892)
         );
  INVX1 U10547 ( .A(n12595), .Y(n12770) );
  NAND3X1 U10548 ( .A(n12901), .B(n12820), .C(n12818), .Y(n12595) );
  INVX1 U10549 ( .A(n12759), .Y(n12818) );
  INVX1 U10550 ( .A(n12593), .Y(n12780) );
  NAND2X1 U10551 ( .A(n12902), .B(n12606), .Y(n12593) );
  OAI21X1 U10552 ( .A(n12468), .B(n12903), .C(n12904), .Y(n5133) );
  NAND2X1 U10553 ( .A(N2513), .B(n12905), .Y(n12904) );
  OAI21X1 U10554 ( .A(n12468), .B(n12906), .C(n12907), .Y(n5132) );
  NAND2X1 U10555 ( .A(N2514), .B(n12905), .Y(n12907) );
  OAI21X1 U10556 ( .A(n12468), .B(n12908), .C(n12909), .Y(n5131) );
  NAND2X1 U10557 ( .A(N2515), .B(n12905), .Y(n12909) );
  OAI21X1 U10558 ( .A(n12468), .B(n12910), .C(n12911), .Y(n5130) );
  NAND2X1 U10559 ( .A(N2516), .B(n12905), .Y(n12911) );
  OAI21X1 U10560 ( .A(n12468), .B(n12912), .C(n12913), .Y(n5129) );
  NAND2X1 U10561 ( .A(N2517), .B(n12905), .Y(n12913) );
  OAI21X1 U10562 ( .A(n12468), .B(n12914), .C(n12915), .Y(n5128) );
  NAND2X1 U10563 ( .A(N2518), .B(n12905), .Y(n12915) );
  OAI21X1 U10564 ( .A(n12468), .B(n12916), .C(n12917), .Y(n5127) );
  NAND2X1 U10565 ( .A(N2519), .B(n12905), .Y(n12917) );
  OAI21X1 U10566 ( .A(n12468), .B(n12918), .C(n12919), .Y(n5126) );
  NAND2X1 U10567 ( .A(N2520), .B(n12905), .Y(n12919) );
  OAI21X1 U10568 ( .A(n12468), .B(n12920), .C(n12921), .Y(n5125) );
  NAND2X1 U10569 ( .A(N2521), .B(n12905), .Y(n12921) );
  OAI21X1 U10570 ( .A(n12468), .B(n12922), .C(n12923), .Y(n5124) );
  NAND2X1 U10571 ( .A(N2522), .B(n12905), .Y(n12923) );
  OAI21X1 U10572 ( .A(n12468), .B(n12924), .C(n12925), .Y(n5123) );
  NAND2X1 U10573 ( .A(N2523), .B(n12905), .Y(n12925) );
  OAI21X1 U10574 ( .A(n12468), .B(n12926), .C(n12927), .Y(n5122) );
  NAND2X1 U10575 ( .A(N2524), .B(n12905), .Y(n12927) );
  INVX1 U10576 ( .A(Gy[11]), .Y(n12926) );
  OAI21X1 U10577 ( .A(n12468), .B(n12928), .C(n12929), .Y(n5121) );
  NAND2X1 U10578 ( .A(N2525), .B(n12905), .Y(n12929) );
  INVX1 U10579 ( .A(Gy[12]), .Y(n12928) );
  OAI21X1 U10580 ( .A(n12468), .B(n12930), .C(n12931), .Y(n5120) );
  NAND2X1 U10581 ( .A(N2526), .B(n12905), .Y(n12931) );
  INVX1 U10582 ( .A(Gy[13]), .Y(n12930) );
  OAI21X1 U10583 ( .A(n12468), .B(n12932), .C(n12933), .Y(n5119) );
  NAND2X1 U10584 ( .A(N2527), .B(n12905), .Y(n12933) );
  INVX1 U10585 ( .A(Gy[14]), .Y(n12932) );
  OAI21X1 U10586 ( .A(n12468), .B(n12934), .C(n12935), .Y(n5118) );
  NAND2X1 U10587 ( .A(N2528), .B(n12905), .Y(n12935) );
  INVX1 U10588 ( .A(Gy[15]), .Y(n12934) );
  OAI21X1 U10589 ( .A(n12468), .B(n12936), .C(n12937), .Y(n5117) );
  NAND2X1 U10590 ( .A(N2529), .B(n12905), .Y(n12937) );
  INVX1 U10591 ( .A(Gy[16]), .Y(n12936) );
  OAI21X1 U10592 ( .A(n12468), .B(n12938), .C(n12939), .Y(n5116) );
  NAND2X1 U10593 ( .A(N2530), .B(n12905), .Y(n12939) );
  INVX1 U10594 ( .A(Gy[17]), .Y(n12938) );
  OAI21X1 U10595 ( .A(n12468), .B(n12940), .C(n12941), .Y(n5115) );
  NAND2X1 U10596 ( .A(N2531), .B(n12905), .Y(n12941) );
  INVX1 U10597 ( .A(Gy[18]), .Y(n12940) );
  OAI21X1 U10598 ( .A(n12468), .B(n12942), .C(n12943), .Y(n5114) );
  NAND2X1 U10599 ( .A(N2532), .B(n12905), .Y(n12943) );
  INVX1 U10600 ( .A(Gy[19]), .Y(n12942) );
  OAI21X1 U10601 ( .A(n12468), .B(n12944), .C(n12945), .Y(n5113) );
  NAND2X1 U10602 ( .A(N2533), .B(n12905), .Y(n12945) );
  INVX1 U10603 ( .A(Gy[20]), .Y(n12944) );
  OAI21X1 U10604 ( .A(n12468), .B(n12946), .C(n12947), .Y(n5112) );
  NAND2X1 U10605 ( .A(N2534), .B(n12905), .Y(n12947) );
  INVX1 U10606 ( .A(Gy[21]), .Y(n12946) );
  OAI21X1 U10607 ( .A(n12468), .B(n12948), .C(n12949), .Y(n5111) );
  NAND2X1 U10608 ( .A(N2535), .B(n12905), .Y(n12949) );
  INVX1 U10609 ( .A(Gy[22]), .Y(n12948) );
  OAI21X1 U10610 ( .A(n12468), .B(n12950), .C(n12951), .Y(n5110) );
  NAND2X1 U10611 ( .A(N2536), .B(n12905), .Y(n12951) );
  INVX1 U10612 ( .A(Gy[23]), .Y(n12950) );
  OAI21X1 U10613 ( .A(n12468), .B(n12952), .C(n12953), .Y(n5109) );
  NAND2X1 U10614 ( .A(N2537), .B(n12905), .Y(n12953) );
  INVX1 U10615 ( .A(Gy[24]), .Y(n12952) );
  OAI21X1 U10616 ( .A(n12468), .B(n12954), .C(n12955), .Y(n5108) );
  NAND2X1 U10617 ( .A(N2538), .B(n12905), .Y(n12955) );
  INVX1 U10618 ( .A(Gy[25]), .Y(n12954) );
  OAI21X1 U10619 ( .A(n12468), .B(n12956), .C(n12957), .Y(n5107) );
  NAND2X1 U10620 ( .A(N2539), .B(n12905), .Y(n12957) );
  INVX1 U10621 ( .A(Gy[26]), .Y(n12956) );
  OAI21X1 U10622 ( .A(n12468), .B(n12958), .C(n12959), .Y(n5106) );
  NAND2X1 U10623 ( .A(N2540), .B(n12905), .Y(n12959) );
  INVX1 U10624 ( .A(Gy[27]), .Y(n12958) );
  OAI21X1 U10625 ( .A(n12468), .B(n12960), .C(n12961), .Y(n5105) );
  NAND2X1 U10626 ( .A(N2541), .B(n12905), .Y(n12961) );
  INVX1 U10627 ( .A(Gy[28]), .Y(n12960) );
  OAI21X1 U10628 ( .A(n12468), .B(n12962), .C(n12963), .Y(n5104) );
  NAND2X1 U10629 ( .A(N2542), .B(n12905), .Y(n12963) );
  INVX1 U10630 ( .A(Gy[29]), .Y(n12962) );
  OAI21X1 U10631 ( .A(n12468), .B(n12964), .C(n12965), .Y(n5103) );
  NAND2X1 U10632 ( .A(N2543), .B(n12905), .Y(n12965) );
  INVX1 U10633 ( .A(Gy[30]), .Y(n12964) );
  OAI21X1 U10634 ( .A(n12468), .B(n12966), .C(n12967), .Y(n5102) );
  NAND2X1 U10635 ( .A(N2544), .B(n12905), .Y(n12967) );
  INVX1 U10636 ( .A(Gy[31]), .Y(n12966) );
  OAI21X1 U10637 ( .A(n15430), .B(n12968), .C(n12969), .Y(n5101) );
  INVX1 U10638 ( .A(N4418), .Y(n15430) );
  OAI21X1 U10639 ( .A(n15431), .B(n12968), .C(n12969), .Y(n5100) );
  INVX1 U10640 ( .A(N4415), .Y(n15431) );
  OAI21X1 U10641 ( .A(n15432), .B(n12968), .C(n12969), .Y(n5099) );
  INVX1 U10642 ( .A(N4412), .Y(n15432) );
  OAI21X1 U10643 ( .A(n15433), .B(n12968), .C(n12969), .Y(n5098) );
  INVX1 U10644 ( .A(N4409), .Y(n15433) );
  OAI21X1 U10645 ( .A(n15434), .B(n12968), .C(n12969), .Y(n5097) );
  INVX1 U10646 ( .A(N4406), .Y(n15434) );
  OAI21X1 U10647 ( .A(n15435), .B(n12968), .C(n12969), .Y(n5096) );
  INVX1 U10648 ( .A(N4403), .Y(n15435) );
  OAI21X1 U10649 ( .A(n15436), .B(n12968), .C(n12969), .Y(n5095) );
  INVX1 U10650 ( .A(N4400), .Y(n15436) );
  OAI21X1 U10651 ( .A(n15437), .B(n12968), .C(n12969), .Y(n5094) );
  NAND2X1 U10652 ( .A(n12968), .B(n12477), .Y(n12969) );
  INVX1 U10653 ( .A(N4397), .Y(n15437) );
  OAI21X1 U10654 ( .A(n12473), .B(n12970), .C(n12971), .Y(n5093) );
  AOI22X1 U10655 ( .A(N2308), .B(n12972), .C(Gx[8]), .D(n12973), .Y(n12971) );
  OAI21X1 U10656 ( .A(n15438), .B(n12473), .C(n12974), .Y(n5092) );
  AOI22X1 U10657 ( .A(N2648), .B(n12975), .C(n12976), .D(Gy[0]), .Y(n12974) );
  INVX1 U10658 ( .A(N4465), .Y(n15438) );
  OAI21X1 U10659 ( .A(n15439), .B(n12473), .C(n12977), .Y(n5091) );
  AOI22X1 U10660 ( .A(N2746), .B(n12975), .C(n12976), .D(Gy[1]), .Y(n12977) );
  INVX1 U10661 ( .A(N4462), .Y(n15439) );
  OAI21X1 U10662 ( .A(n15440), .B(n12473), .C(n12978), .Y(n5090) );
  AOI22X1 U10663 ( .A(N2747), .B(n12975), .C(n12976), .D(Gy[2]), .Y(n12978) );
  INVX1 U10664 ( .A(N4459), .Y(n15440) );
  OAI21X1 U10665 ( .A(n15441), .B(n12473), .C(n12979), .Y(n5089) );
  AOI22X1 U10666 ( .A(N2748), .B(n12975), .C(n12976), .D(Gy[3]), .Y(n12979) );
  INVX1 U10667 ( .A(N4456), .Y(n15441) );
  OAI21X1 U10668 ( .A(n15442), .B(n12473), .C(n12980), .Y(n5088) );
  AOI22X1 U10669 ( .A(N2749), .B(n12975), .C(n12976), .D(Gy[4]), .Y(n12980) );
  INVX1 U10670 ( .A(N4453), .Y(n15442) );
  OAI21X1 U10671 ( .A(n15443), .B(n12473), .C(n12981), .Y(n5087) );
  AOI22X1 U10672 ( .A(n12975), .B(N2750), .C(n12976), .D(Gy[5]), .Y(n12981) );
  INVX1 U10673 ( .A(N4450), .Y(n15443) );
  OAI21X1 U10674 ( .A(n15444), .B(n12473), .C(n12982), .Y(n5086) );
  AOI22X1 U10675 ( .A(n12975), .B(N2751), .C(n12976), .D(Gy[6]), .Y(n12982) );
  INVX1 U10676 ( .A(N4447), .Y(n15444) );
  OAI21X1 U10677 ( .A(n15445), .B(n12473), .C(n12983), .Y(n5085) );
  AOI22X1 U10678 ( .A(n12975), .B(N2752), .C(n12976), .D(Gy[7]), .Y(n12983) );
  INVX1 U10679 ( .A(N4444), .Y(n15445) );
  OAI21X1 U10680 ( .A(n12984), .B(n12473), .C(n12985), .Y(n5084) );
  AOI22X1 U10681 ( .A(n12972), .B(N2753), .C(n12973), .D(Gy[8]), .Y(n12985) );
  OAI21X1 U10682 ( .A(n12986), .B(n12473), .C(n12987), .Y(n5083) );
  AOI22X1 U10683 ( .A(N2754), .B(n12972), .C(n12973), .D(Gy[9]), .Y(n12987) );
  OAI21X1 U10684 ( .A(n12988), .B(n12473), .C(n12989), .Y(n5082) );
  AOI22X1 U10685 ( .A(N2755), .B(n12972), .C(n12973), .D(Gy[10]), .Y(n12989)
         );
  OAI21X1 U10686 ( .A(n12990), .B(n12473), .C(n12991), .Y(n5081) );
  AOI22X1 U10687 ( .A(N2756), .B(n12972), .C(n12973), .D(Gy[11]), .Y(n12991)
         );
  OAI21X1 U10688 ( .A(n12992), .B(n12473), .C(n12993), .Y(n5080) );
  AOI22X1 U10689 ( .A(N2757), .B(n12972), .C(n12973), .D(Gy[12]), .Y(n12993)
         );
  OAI21X1 U10690 ( .A(n12994), .B(n12473), .C(n12995), .Y(n5079) );
  AOI22X1 U10691 ( .A(N2758), .B(n12972), .C(n12973), .D(Gy[13]), .Y(n12995)
         );
  OAI21X1 U10692 ( .A(n12996), .B(n12473), .C(n12997), .Y(n5078) );
  AOI22X1 U10693 ( .A(N2759), .B(n12972), .C(n12973), .D(Gy[14]), .Y(n12997)
         );
  OAI21X1 U10694 ( .A(n12998), .B(n12473), .C(n12999), .Y(n5077) );
  AOI22X1 U10695 ( .A(N2760), .B(n12972), .C(n12973), .D(Gy[15]), .Y(n12999)
         );
  OAI21X1 U10696 ( .A(n13000), .B(n12473), .C(n13001), .Y(n5076) );
  AOI22X1 U10697 ( .A(N2761), .B(n12972), .C(n12973), .D(Gy[16]), .Y(n13001)
         );
  OAI21X1 U10698 ( .A(n13002), .B(n12473), .C(n13003), .Y(n5075) );
  AOI22X1 U10699 ( .A(N2762), .B(n12972), .C(n12973), .D(Gy[17]), .Y(n13003)
         );
  OAI21X1 U10700 ( .A(n13004), .B(n12473), .C(n13005), .Y(n5074) );
  AOI22X1 U10701 ( .A(N2763), .B(n12972), .C(n12973), .D(Gy[18]), .Y(n13005)
         );
  OAI21X1 U10702 ( .A(n13006), .B(n12473), .C(n13007), .Y(n5073) );
  AOI22X1 U10703 ( .A(N2764), .B(n12972), .C(n12973), .D(Gy[19]), .Y(n13007)
         );
  OAI21X1 U10704 ( .A(n13008), .B(n12473), .C(n13009), .Y(n5072) );
  AOI22X1 U10705 ( .A(N2765), .B(n12972), .C(n12973), .D(Gy[20]), .Y(n13009)
         );
  OAI21X1 U10706 ( .A(n13010), .B(n12473), .C(n13011), .Y(n5071) );
  AOI22X1 U10707 ( .A(N2766), .B(n12972), .C(n12973), .D(Gy[21]), .Y(n13011)
         );
  OAI21X1 U10708 ( .A(n13012), .B(n12473), .C(n13013), .Y(n5070) );
  AOI22X1 U10709 ( .A(N2767), .B(n12972), .C(n12973), .D(Gy[22]), .Y(n13013)
         );
  OAI21X1 U10710 ( .A(n13014), .B(n12473), .C(n13015), .Y(n5069) );
  AOI22X1 U10711 ( .A(N2768), .B(n12972), .C(n12973), .D(Gy[23]), .Y(n13015)
         );
  OAI21X1 U10712 ( .A(n13016), .B(n12473), .C(n13017), .Y(n5068) );
  AOI22X1 U10713 ( .A(N2769), .B(n12972), .C(n12973), .D(Gy[24]), .Y(n13017)
         );
  OAI21X1 U10714 ( .A(n13018), .B(n12473), .C(n13019), .Y(n5067) );
  AOI22X1 U10715 ( .A(N2770), .B(n12972), .C(n12973), .D(Gy[25]), .Y(n13019)
         );
  OAI21X1 U10716 ( .A(n13020), .B(n12473), .C(n13021), .Y(n5066) );
  AOI22X1 U10717 ( .A(N2771), .B(n12972), .C(n12973), .D(Gy[26]), .Y(n13021)
         );
  OAI21X1 U10718 ( .A(n13022), .B(n12473), .C(n13023), .Y(n5065) );
  AOI22X1 U10719 ( .A(N2772), .B(n12972), .C(n12973), .D(Gy[27]), .Y(n13023)
         );
  OAI21X1 U10720 ( .A(n13024), .B(n12473), .C(n13025), .Y(n5064) );
  AOI22X1 U10721 ( .A(N2773), .B(n12972), .C(n12973), .D(Gy[28]), .Y(n13025)
         );
  OAI21X1 U10722 ( .A(n13026), .B(n12473), .C(n13027), .Y(n5063) );
  AOI22X1 U10723 ( .A(N2774), .B(n12972), .C(n12973), .D(Gy[29]), .Y(n13027)
         );
  OAI21X1 U10724 ( .A(n13028), .B(n12473), .C(n13029), .Y(n5062) );
  AOI22X1 U10725 ( .A(N2775), .B(n12972), .C(n12973), .D(Gy[30]), .Y(n13029)
         );
  OAI22X1 U10726 ( .A(n13030), .B(n12473), .C(n13031), .D(n13032), .Y(n5061)
         );
  OAI22X1 U10727 ( .A(n12468), .B(n13033), .C(n13034), .D(n13035), .Y(n5060)
         );
  INVX1 U10728 ( .A(N2300), .Y(n13035) );
  OAI21X1 U10729 ( .A(n15446), .B(n12473), .C(n13036), .Y(n5059) );
  AOI22X1 U10730 ( .A(N2300), .B(n12975), .C(Gx[0]), .D(n12976), .Y(n13036) );
  INVX1 U10731 ( .A(N4393), .Y(n15446) );
  OAI22X1 U10732 ( .A(n12468), .B(n13037), .C(n13034), .D(n13038), .Y(n5058)
         );
  INVX1 U10733 ( .A(N2301), .Y(n13038) );
  OAI21X1 U10734 ( .A(n15447), .B(n12473), .C(n13039), .Y(n5057) );
  AOI22X1 U10735 ( .A(N2301), .B(n12975), .C(Gx[1]), .D(n12976), .Y(n13039) );
  INVX1 U10736 ( .A(N4390), .Y(n15447) );
  OAI22X1 U10737 ( .A(n12468), .B(n13040), .C(n13034), .D(n13041), .Y(n5056)
         );
  INVX1 U10738 ( .A(N2302), .Y(n13041) );
  OAI21X1 U10739 ( .A(n15448), .B(n12473), .C(n13042), .Y(n5055) );
  AOI22X1 U10740 ( .A(N2302), .B(n12975), .C(Gx[2]), .D(n12976), .Y(n13042) );
  INVX1 U10741 ( .A(N4387), .Y(n15448) );
  OAI22X1 U10742 ( .A(n12468), .B(n13043), .C(n13034), .D(n13044), .Y(n5054)
         );
  INVX1 U10743 ( .A(N2303), .Y(n13044) );
  OAI21X1 U10744 ( .A(n15449), .B(n12473), .C(n13045), .Y(n5053) );
  AOI22X1 U10745 ( .A(N2303), .B(n12975), .C(Gx[3]), .D(n12976), .Y(n13045) );
  INVX1 U10746 ( .A(N4384), .Y(n15449) );
  OAI22X1 U10747 ( .A(n12468), .B(n13046), .C(n13034), .D(n13047), .Y(n5052)
         );
  INVX1 U10748 ( .A(N2304), .Y(n13047) );
  OAI21X1 U10749 ( .A(n15450), .B(n12473), .C(n13048), .Y(n5051) );
  AOI22X1 U10750 ( .A(N2304), .B(n12975), .C(Gx[4]), .D(n12976), .Y(n13048) );
  INVX1 U10751 ( .A(N4381), .Y(n15450) );
  OAI22X1 U10752 ( .A(n12468), .B(n13049), .C(n13034), .D(n13050), .Y(n5050)
         );
  INVX1 U10753 ( .A(N2305), .Y(n13050) );
  OAI21X1 U10754 ( .A(n15451), .B(n12473), .C(n13051), .Y(n5049) );
  AOI22X1 U10755 ( .A(N2305), .B(n12975), .C(Gx[5]), .D(n12976), .Y(n13051) );
  INVX1 U10756 ( .A(N4378), .Y(n15451) );
  OAI22X1 U10757 ( .A(n12468), .B(n13052), .C(n13034), .D(n13053), .Y(n5048)
         );
  INVX1 U10758 ( .A(N2306), .Y(n13053) );
  OAI21X1 U10759 ( .A(n15452), .B(n12473), .C(n13054), .Y(n5047) );
  AOI22X1 U10760 ( .A(N2306), .B(n12975), .C(Gx[6]), .D(n12976), .Y(n13054) );
  INVX1 U10761 ( .A(N4375), .Y(n15452) );
  OAI22X1 U10762 ( .A(n12468), .B(n13055), .C(n13034), .D(n13056), .Y(n5046)
         );
  INVX1 U10763 ( .A(N2307), .Y(n13056) );
  OAI21X1 U10764 ( .A(n15453), .B(n12473), .C(n13057), .Y(n5045) );
  AOI22X1 U10765 ( .A(N2307), .B(n12975), .C(Gx[7]), .D(n12976), .Y(n13057) );
  AND2X1 U10766 ( .A(n12473), .B(n13058), .Y(n12975) );
  INVX1 U10767 ( .A(N4372), .Y(n15453) );
  OAI22X1 U10768 ( .A(n12468), .B(n13059), .C(n13034), .D(n13060), .Y(n5044)
         );
  INVX1 U10769 ( .A(N2308), .Y(n13060) );
  OAI22X1 U10770 ( .A(n12468), .B(n13061), .C(n13034), .D(n13062), .Y(n5043)
         );
  INVX1 U10771 ( .A(N2309), .Y(n13062) );
  OAI21X1 U10772 ( .A(n12473), .B(n13063), .C(n13064), .Y(n5042) );
  AOI22X1 U10773 ( .A(N2309), .B(n12972), .C(Gx[9]), .D(n12973), .Y(n13064) );
  OAI22X1 U10774 ( .A(n12468), .B(n13065), .C(n13034), .D(n13066), .Y(n5041)
         );
  INVX1 U10775 ( .A(N2310), .Y(n13066) );
  OAI21X1 U10776 ( .A(n15454), .B(n12968), .C(n13067), .Y(n5040) );
  AOI22X1 U10777 ( .A(N2561), .B(n13068), .C(N2569), .D(n13069), .Y(n13067) );
  INVX1 U10778 ( .A(N4417), .Y(n15454) );
  OAI21X1 U10779 ( .A(n15455), .B(n12968), .C(n13070), .Y(n5039) );
  AOI22X1 U10780 ( .A(N2562), .B(n13068), .C(N2570), .D(n13069), .Y(n13070) );
  INVX1 U10781 ( .A(N4414), .Y(n15455) );
  OAI21X1 U10782 ( .A(n15456), .B(n12968), .C(n13071), .Y(n5038) );
  AOI22X1 U10783 ( .A(N2563), .B(n13068), .C(N2571), .D(n13069), .Y(n13071) );
  INVX1 U10784 ( .A(N4411), .Y(n15456) );
  OAI21X1 U10785 ( .A(n15457), .B(n12968), .C(n13072), .Y(n5037) );
  AOI22X1 U10786 ( .A(N2564), .B(n13068), .C(N2572), .D(n13069), .Y(n13072) );
  INVX1 U10787 ( .A(N4408), .Y(n15457) );
  OAI21X1 U10788 ( .A(n15458), .B(n12968), .C(n13073), .Y(n5036) );
  AOI22X1 U10789 ( .A(N2565), .B(n13068), .C(N2573), .D(n13069), .Y(n13073) );
  INVX1 U10790 ( .A(N4405), .Y(n15458) );
  OAI21X1 U10791 ( .A(n15459), .B(n12968), .C(n13074), .Y(n5035) );
  AOI22X1 U10792 ( .A(N2566), .B(n13068), .C(N2574), .D(n13069), .Y(n13074) );
  INVX1 U10793 ( .A(N4402), .Y(n15459) );
  OAI21X1 U10794 ( .A(n15460), .B(n12968), .C(n13075), .Y(n5034) );
  AOI22X1 U10795 ( .A(N2567), .B(n13068), .C(N2575), .D(n13069), .Y(n13075) );
  INVX1 U10796 ( .A(N4399), .Y(n15460) );
  OAI21X1 U10797 ( .A(n15461), .B(n12968), .C(n13076), .Y(n5033) );
  AOI22X1 U10798 ( .A(N2568), .B(n13068), .C(N2576), .D(n13069), .Y(n13076) );
  AOI21X1 U10799 ( .A(n13058), .B(n8303), .C(n13077), .Y(n13069) );
  INVX1 U10800 ( .A(n13078), .Y(n13068) );
  NAND3X1 U10801 ( .A(n12968), .B(n13058), .C(N2549), .Y(n13078) );
  INVX1 U10802 ( .A(n13077), .Y(n12968) );
  INVX1 U10803 ( .A(N4396), .Y(n15461) );
  OAI21X1 U10804 ( .A(n12473), .B(n13079), .C(n13080), .Y(n5032) );
  AOI22X1 U10805 ( .A(N2310), .B(n12972), .C(Gx[10]), .D(n12973), .Y(n13080)
         );
  OAI22X1 U10806 ( .A(n12468), .B(n13081), .C(n13034), .D(n13082), .Y(n5031)
         );
  INVX1 U10807 ( .A(N2311), .Y(n13082) );
  OAI21X1 U10808 ( .A(n12473), .B(n13083), .C(n13084), .Y(n5030) );
  AOI22X1 U10809 ( .A(N2311), .B(n12972), .C(Gx[11]), .D(n12973), .Y(n13084)
         );
  OAI22X1 U10810 ( .A(n12468), .B(n13085), .C(n13034), .D(n13086), .Y(n5029)
         );
  INVX1 U10811 ( .A(N2312), .Y(n13086) );
  OAI21X1 U10812 ( .A(n12473), .B(n13087), .C(n13088), .Y(n5028) );
  AOI22X1 U10813 ( .A(N2312), .B(n12972), .C(Gx[12]), .D(n12973), .Y(n13088)
         );
  OAI22X1 U10814 ( .A(n12468), .B(n13089), .C(n13034), .D(n13090), .Y(n5027)
         );
  INVX1 U10815 ( .A(N2313), .Y(n13090) );
  OAI21X1 U10816 ( .A(n12473), .B(n13091), .C(n13092), .Y(n5026) );
  AOI22X1 U10817 ( .A(N2313), .B(n12972), .C(Gx[13]), .D(n12973), .Y(n13092)
         );
  OAI22X1 U10818 ( .A(n12468), .B(n13093), .C(n13034), .D(n13094), .Y(n5025)
         );
  INVX1 U10819 ( .A(N2314), .Y(n13094) );
  OAI21X1 U10820 ( .A(n12473), .B(n13095), .C(n13096), .Y(n5024) );
  AOI22X1 U10821 ( .A(N2314), .B(n12972), .C(Gx[14]), .D(n12973), .Y(n13096)
         );
  OAI22X1 U10822 ( .A(n12468), .B(n13097), .C(n13034), .D(n13098), .Y(n5023)
         );
  INVX1 U10823 ( .A(N2315), .Y(n13098) );
  OAI21X1 U10824 ( .A(n12473), .B(n13099), .C(n13100), .Y(n5022) );
  AOI22X1 U10825 ( .A(N2315), .B(n12972), .C(Gx[15]), .D(n12973), .Y(n13100)
         );
  OAI22X1 U10826 ( .A(n12468), .B(n13101), .C(n13034), .D(n13102), .Y(n5021)
         );
  INVX1 U10827 ( .A(N2316), .Y(n13102) );
  OAI21X1 U10828 ( .A(n12473), .B(n13103), .C(n13104), .Y(n5020) );
  AOI22X1 U10829 ( .A(N2316), .B(n12972), .C(Gx[16]), .D(n12973), .Y(n13104)
         );
  OAI22X1 U10830 ( .A(n12468), .B(n13105), .C(n13034), .D(n13106), .Y(n5019)
         );
  INVX1 U10831 ( .A(N2317), .Y(n13106) );
  OAI21X1 U10832 ( .A(n12473), .B(n13107), .C(n13108), .Y(n5018) );
  AOI22X1 U10833 ( .A(N2317), .B(n12972), .C(Gx[17]), .D(n12973), .Y(n13108)
         );
  OAI22X1 U10834 ( .A(n12468), .B(n13109), .C(n13034), .D(n13110), .Y(n5017)
         );
  INVX1 U10835 ( .A(N2318), .Y(n13110) );
  OAI21X1 U10836 ( .A(n12473), .B(n13111), .C(n13112), .Y(n5016) );
  AOI22X1 U10837 ( .A(N2318), .B(n12972), .C(Gx[18]), .D(n12973), .Y(n13112)
         );
  OAI22X1 U10838 ( .A(n12468), .B(n13113), .C(n13034), .D(n13114), .Y(n5015)
         );
  INVX1 U10839 ( .A(N2319), .Y(n13114) );
  OAI21X1 U10840 ( .A(n12473), .B(n13115), .C(n13116), .Y(n5014) );
  AOI22X1 U10841 ( .A(N2319), .B(n12972), .C(Gx[19]), .D(n12973), .Y(n13116)
         );
  OAI22X1 U10842 ( .A(n12468), .B(n13117), .C(n13034), .D(n13118), .Y(n5013)
         );
  INVX1 U10843 ( .A(N2320), .Y(n13118) );
  OAI21X1 U10844 ( .A(n12473), .B(n13119), .C(n13120), .Y(n5012) );
  AOI22X1 U10845 ( .A(N2320), .B(n12972), .C(Gx[20]), .D(n12973), .Y(n13120)
         );
  OAI22X1 U10846 ( .A(n12468), .B(n13121), .C(n13034), .D(n13122), .Y(n5011)
         );
  INVX1 U10847 ( .A(N2321), .Y(n13122) );
  OAI21X1 U10848 ( .A(n12473), .B(n13123), .C(n13124), .Y(n5010) );
  AOI22X1 U10849 ( .A(N2321), .B(n12972), .C(Gx[21]), .D(n12973), .Y(n13124)
         );
  OAI22X1 U10850 ( .A(n12468), .B(n13125), .C(n13034), .D(n13126), .Y(n5009)
         );
  INVX1 U10851 ( .A(N2322), .Y(n13126) );
  OAI21X1 U10852 ( .A(n12473), .B(n13127), .C(n13128), .Y(n5008) );
  AOI22X1 U10853 ( .A(N2322), .B(n12972), .C(Gx[22]), .D(n12973), .Y(n13128)
         );
  OAI22X1 U10854 ( .A(n12468), .B(n13129), .C(n13034), .D(n13130), .Y(n5007)
         );
  INVX1 U10855 ( .A(N2323), .Y(n13130) );
  OAI21X1 U10856 ( .A(n12473), .B(n13131), .C(n13132), .Y(n5006) );
  AOI22X1 U10857 ( .A(N2323), .B(n12972), .C(Gx[23]), .D(n12973), .Y(n13132)
         );
  OAI22X1 U10858 ( .A(n12468), .B(n13133), .C(n13034), .D(n13134), .Y(n5005)
         );
  INVX1 U10859 ( .A(N2324), .Y(n13134) );
  OAI21X1 U10860 ( .A(n12473), .B(n13135), .C(n13136), .Y(n5004) );
  AOI22X1 U10861 ( .A(N2324), .B(n12972), .C(Gx[24]), .D(n12973), .Y(n13136)
         );
  OAI22X1 U10862 ( .A(n12468), .B(n13137), .C(n13034), .D(n13138), .Y(n5003)
         );
  INVX1 U10863 ( .A(N2325), .Y(n13138) );
  OAI21X1 U10864 ( .A(n12473), .B(n13139), .C(n13140), .Y(n5002) );
  AOI22X1 U10865 ( .A(N2325), .B(n12972), .C(Gx[25]), .D(n12973), .Y(n13140)
         );
  OAI22X1 U10866 ( .A(n12468), .B(n13141), .C(n13034), .D(n13142), .Y(n5001)
         );
  INVX1 U10867 ( .A(N2326), .Y(n13142) );
  OAI21X1 U10868 ( .A(n12473), .B(n13143), .C(n13144), .Y(n5000) );
  AOI22X1 U10869 ( .A(N2326), .B(n12972), .C(Gx[26]), .D(n12973), .Y(n13144)
         );
  OAI22X1 U10870 ( .A(n12468), .B(n13145), .C(n13034), .D(n13146), .Y(n4999)
         );
  INVX1 U10871 ( .A(N2327), .Y(n13146) );
  OAI21X1 U10872 ( .A(n12473), .B(n13147), .C(n13148), .Y(n4998) );
  AOI22X1 U10873 ( .A(N2327), .B(n12972), .C(Gx[27]), .D(n12973), .Y(n13148)
         );
  OAI22X1 U10874 ( .A(n12468), .B(n13149), .C(n13034), .D(n13150), .Y(n4997)
         );
  INVX1 U10875 ( .A(N2328), .Y(n13150) );
  OAI21X1 U10876 ( .A(n12473), .B(n13151), .C(n13152), .Y(n4996) );
  AOI22X1 U10877 ( .A(N2328), .B(n12972), .C(Gx[28]), .D(n12973), .Y(n13152)
         );
  OAI22X1 U10878 ( .A(n12468), .B(n13153), .C(n13034), .D(n13154), .Y(n4995)
         );
  INVX1 U10879 ( .A(N2329), .Y(n13154) );
  OAI21X1 U10880 ( .A(n12473), .B(n13155), .C(n13156), .Y(n4994) );
  AOI22X1 U10881 ( .A(N2329), .B(n12972), .C(Gx[29]), .D(n12973), .Y(n13156)
         );
  OAI22X1 U10882 ( .A(n12468), .B(n13157), .C(n13034), .D(n13158), .Y(n4993)
         );
  INVX1 U10883 ( .A(N2330), .Y(n13158) );
  OAI21X1 U10884 ( .A(n12473), .B(n13159), .C(n13160), .Y(n4992) );
  AOI22X1 U10885 ( .A(N2330), .B(n12972), .C(Gx[30]), .D(n12973), .Y(n13160)
         );
  OAI22X1 U10886 ( .A(n12468), .B(n13161), .C(n13034), .D(n13162), .Y(n4991)
         );
  INVX1 U10887 ( .A(N2331), .Y(n13162) );
  NOR2X1 U10888 ( .A(n13077), .B(n12462), .Y(n12905) );
  OAI21X1 U10889 ( .A(n13163), .B(n12473), .C(n13164), .Y(n4990) );
  AOI22X1 U10890 ( .A(N2331), .B(n12972), .C(Gx[31]), .D(n12973), .Y(n13164)
         );
  NAND2X1 U10891 ( .A(n12475), .B(n12473), .Y(n13031) );
  OAI21X1 U10892 ( .A(n12680), .B(n12568), .C(n13077), .Y(n12571) );
  NAND3X1 U10893 ( .A(n13166), .B(n12573), .C(n12668), .Y(n13077) );
  MUX2X1 U10894 ( .B(n12577), .A(n12555), .S(n13167), .Y(n4989) );
  MUX2X1 U10895 ( .B(n12580), .A(n13168), .S(n13167), .Y(n4988) );
  MUX2X1 U10896 ( .B(n12582), .A(n13169), .S(n13167), .Y(n4987) );
  MUX2X1 U10897 ( .B(n12584), .A(n13170), .S(n13167), .Y(n4986) );
  MUX2X1 U10898 ( .B(n12586), .A(n13171), .S(n13167), .Y(n4985) );
  MUX2X1 U10899 ( .B(n12588), .A(n13172), .S(n13167), .Y(n4984) );
  MUX2X1 U10900 ( .B(n12590), .A(n13173), .S(n13167), .Y(n4983) );
  MUX2X1 U10901 ( .B(n12592), .A(n13174), .S(n13167), .Y(n4982) );
  AOI22X1 U10902 ( .A(n12802), .B(n13175), .C(n12711), .D(n12792), .Y(n13167)
         );
  MUX2X1 U10903 ( .B(n12577), .A(n13176), .S(n13177), .Y(n4981) );
  NAND2X1 U10904 ( .A(InData[0]), .B(n12494), .Y(n12577) );
  MUX2X1 U10905 ( .B(n12580), .A(n13178), .S(n13177), .Y(n4980) );
  NAND2X1 U10906 ( .A(InData[1]), .B(n12494), .Y(n12580) );
  MUX2X1 U10907 ( .B(n12582), .A(n13179), .S(n13177), .Y(n4979) );
  NAND2X1 U10908 ( .A(InData[2]), .B(n12494), .Y(n12582) );
  MUX2X1 U10909 ( .B(n12584), .A(n13180), .S(n13177), .Y(n4978) );
  NAND2X1 U10910 ( .A(InData[3]), .B(n12494), .Y(n12584) );
  MUX2X1 U10911 ( .B(n12586), .A(n13181), .S(n13177), .Y(n4977) );
  NAND2X1 U10912 ( .A(InData[4]), .B(n12494), .Y(n12586) );
  MUX2X1 U10913 ( .B(n12588), .A(n13182), .S(n13177), .Y(n4976) );
  NAND2X1 U10914 ( .A(InData[5]), .B(n12494), .Y(n12588) );
  MUX2X1 U10915 ( .B(n12590), .A(n13183), .S(n13177), .Y(n4975) );
  NAND2X1 U10916 ( .A(InData[6]), .B(n12494), .Y(n12590) );
  MUX2X1 U10917 ( .B(n12592), .A(n13184), .S(n13177), .Y(n4974) );
  AOI22X1 U10918 ( .A(n12802), .B(n13185), .C(n12722), .D(n12792), .Y(n13177)
         );
  NOR3X1 U10919 ( .A(n12759), .B(n12901), .C(n12820), .Y(n12792) );
  NAND3X1 U10920 ( .A(n12668), .B(n12689), .C(n15327), .Y(n12759) );
  XOR2X1 U10921 ( .A(N3194), .B(n13186), .Y(n12689) );
  NOR2X1 U10922 ( .A(n13187), .B(n13188), .Y(n13186) );
  AND2X1 U10923 ( .A(n13189), .B(n12606), .Y(n12802) );
  OAI21X1 U10924 ( .A(n12684), .B(n13190), .C(n12679), .Y(n12606) );
  NAND3X1 U10925 ( .A(n13191), .B(n13192), .C(n13193), .Y(n12679) );
  NAND2X1 U10926 ( .A(n15327), .B(n12668), .Y(n13190) );
  NAND2X1 U10927 ( .A(n13194), .B(n13195), .Y(n12684) );
  NAND2X1 U10928 ( .A(InData[7]), .B(n12494), .Y(n12592) );
  OAI21X1 U10929 ( .A(n15462), .B(n13196), .C(n13197), .Y(n4973) );
  INVX1 U10930 ( .A(N4441), .Y(n15462) );
  OAI21X1 U10931 ( .A(n15463), .B(n13196), .C(n13198), .Y(n4972) );
  INVX1 U10932 ( .A(N4442), .Y(n15463) );
  NAND2X1 U10933 ( .A(n13199), .B(n13200), .Y(n4971) );
  MUX2X1 U10934 ( .B(N4438), .A(n13201), .S(n13196), .Y(n13199) );
  OAI21X1 U10935 ( .A(n13202), .B(n13203), .C(n13204), .Y(n13201) );
  INVX1 U10936 ( .A(N2874), .Y(n13203) );
  OAI21X1 U10937 ( .A(n15465), .B(n13196), .C(n13198), .Y(n4970) );
  INVX1 U10938 ( .A(N4439), .Y(n15465) );
  OAI21X1 U10939 ( .A(n15466), .B(n13196), .C(n13197), .Y(n4969) );
  NOR2X1 U10940 ( .A(n13205), .B(n13206), .Y(n13197) );
  INVX1 U10941 ( .A(n13200), .Y(n13206) );
  INVX1 U10942 ( .A(n13207), .Y(n13205) );
  INVX1 U10943 ( .A(N4435), .Y(n15466) );
  OAI21X1 U10944 ( .A(n15467), .B(n13196), .C(n13198), .Y(n4968) );
  INVX1 U10945 ( .A(N4436), .Y(n15467) );
  OAI21X1 U10946 ( .A(n15469), .B(n13196), .C(n13198), .Y(n4966) );
  INVX1 U10947 ( .A(N4433), .Y(n15469) );
  OAI21X1 U10948 ( .A(n15470), .B(n13196), .C(n13208), .Y(n4965) );
  INVX1 U10949 ( .A(N4429), .Y(n15470) );
  OAI21X1 U10950 ( .A(n15471), .B(n13196), .C(n13198), .Y(n4964) );
  INVX1 U10951 ( .A(N4430), .Y(n15471) );
  OAI21X1 U10952 ( .A(n15472), .B(n13196), .C(n13207), .Y(n4963) );
  NAND3X1 U10953 ( .A(n13209), .B(n12687), .C(n13196), .Y(n13207) );
  INVX1 U10954 ( .A(N4426), .Y(n15472) );
  OAI21X1 U10955 ( .A(n15473), .B(n13196), .C(n13198), .Y(n4962) );
  INVX1 U10956 ( .A(N4427), .Y(n15473) );
  OAI21X1 U10957 ( .A(n15474), .B(n13196), .C(n13208), .Y(n4961) );
  OAI21X1 U10958 ( .A(n13210), .B(n13211), .C(n13196), .Y(n13208) );
  INVX1 U10959 ( .A(n13212), .Y(n13211) );
  INVX1 U10960 ( .A(n13204), .Y(n13210) );
  NAND3X1 U10961 ( .A(N2880), .B(n13213), .C(N2945), .Y(n13204) );
  INVX1 U10962 ( .A(N4423), .Y(n15474) );
  OAI21X1 U10963 ( .A(n15475), .B(n13196), .C(n13198), .Y(n4960) );
  INVX1 U10964 ( .A(N4424), .Y(n15475) );
  OAI21X1 U10965 ( .A(n15476), .B(n13196), .C(n13200), .Y(n4959) );
  NAND3X1 U10966 ( .A(n13214), .B(n13215), .C(n13196), .Y(n13200) );
  INVX1 U10967 ( .A(n13216), .Y(n13214) );
  INVX1 U10968 ( .A(N4420), .Y(n15476) );
  OAI21X1 U10969 ( .A(n15477), .B(n13196), .C(n13198), .Y(n4958) );
  NAND2X1 U10970 ( .A(n13196), .B(n12573), .Y(n13198) );
  INVX1 U10971 ( .A(n13217), .Y(n12573) );
  INVX1 U10972 ( .A(N4421), .Y(n15477) );
  MUX2X1 U10973 ( .B(n15478), .A(n12621), .S(n13218), .Y(n4957) );
  INVX1 U10974 ( .A(N3865), .Y(n15478) );
  OAI21X1 U10975 ( .A(n15479), .B(n13218), .C(n13219), .Y(n4956) );
  INVX1 U10976 ( .A(N3866), .Y(n15479) );
  MUX2X1 U10977 ( .B(n15480), .A(n12631), .S(n13218), .Y(n4955) );
  INVX1 U10978 ( .A(N3862), .Y(n15480) );
  OAI21X1 U10979 ( .A(n15481), .B(n13218), .C(n13219), .Y(n4954) );
  INVX1 U10980 ( .A(N3863), .Y(n15481) );
  MUX2X1 U10981 ( .B(n15482), .A(n12629), .S(n13218), .Y(n4953) );
  INVX1 U10982 ( .A(N3859), .Y(n15482) );
  OAI21X1 U10983 ( .A(n15483), .B(n13218), .C(n13219), .Y(n4952) );
  INVX1 U10984 ( .A(N3860), .Y(n15483) );
  MUX2X1 U10985 ( .B(n15484), .A(n12628), .S(n13218), .Y(n4951) );
  INVX1 U10986 ( .A(N3856), .Y(n15484) );
  OAI21X1 U10987 ( .A(n15485), .B(n13218), .C(n13219), .Y(n4950) );
  INVX1 U10988 ( .A(N3857), .Y(n15485) );
  MUX2X1 U10989 ( .B(n15486), .A(n12627), .S(n13218), .Y(n4949) );
  INVX1 U10990 ( .A(N3853), .Y(n15486) );
  OAI21X1 U10991 ( .A(n15487), .B(n13218), .C(n13219), .Y(n4948) );
  INVX1 U10992 ( .A(N3854), .Y(n15487) );
  MUX2X1 U10993 ( .B(n15488), .A(n12626), .S(n13218), .Y(n4947) );
  INVX1 U10994 ( .A(N3850), .Y(n15488) );
  OAI21X1 U10995 ( .A(n15489), .B(n13218), .C(n13219), .Y(n4946) );
  INVX1 U10996 ( .A(N3851), .Y(n15489) );
  MUX2X1 U10997 ( .B(n15490), .A(n12625), .S(n13218), .Y(n4945) );
  INVX1 U10998 ( .A(N3847), .Y(n15490) );
  OAI21X1 U10999 ( .A(n15491), .B(n13218), .C(n13219), .Y(n4944) );
  INVX1 U11000 ( .A(N3848), .Y(n15491) );
  MUX2X1 U11001 ( .B(n15492), .A(n12624), .S(n13218), .Y(n4943) );
  INVX1 U11002 ( .A(N3844), .Y(n15492) );
  OAI21X1 U11003 ( .A(n15493), .B(n13218), .C(n13219), .Y(n4942) );
  NAND2X1 U11004 ( .A(n13218), .B(n12630), .Y(n13219) );
  NOR2X1 U11005 ( .A(n12723), .B(n13220), .Y(n13218) );
  INVX1 U11006 ( .A(N3845), .Y(n15493) );
  MUX2X1 U11007 ( .B(n15494), .A(n12621), .S(n13221), .Y(n4941) );
  INVX1 U11008 ( .A(N3889), .Y(n15494) );
  OAI21X1 U11009 ( .A(n15495), .B(n13221), .C(n13222), .Y(n4940) );
  INVX1 U11010 ( .A(N3890), .Y(n15495) );
  MUX2X1 U11011 ( .B(n15496), .A(n12631), .S(n13221), .Y(n4939) );
  INVX1 U11012 ( .A(N3886), .Y(n15496) );
  OAI21X1 U11013 ( .A(n15497), .B(n13221), .C(n13222), .Y(n4938) );
  INVX1 U11014 ( .A(N3887), .Y(n15497) );
  MUX2X1 U11015 ( .B(n15498), .A(n12629), .S(n13221), .Y(n4937) );
  INVX1 U11016 ( .A(N3883), .Y(n15498) );
  OAI21X1 U11017 ( .A(n15499), .B(n13221), .C(n13222), .Y(n4936) );
  INVX1 U11018 ( .A(N3884), .Y(n15499) );
  MUX2X1 U11019 ( .B(n15500), .A(n12628), .S(n13221), .Y(n4935) );
  INVX1 U11020 ( .A(N3880), .Y(n15500) );
  OAI21X1 U11021 ( .A(n15501), .B(n13221), .C(n13222), .Y(n4934) );
  INVX1 U11022 ( .A(N3881), .Y(n15501) );
  MUX2X1 U11023 ( .B(n15502), .A(n12627), .S(n13221), .Y(n4933) );
  INVX1 U11024 ( .A(N3877), .Y(n15502) );
  OAI21X1 U11025 ( .A(n15503), .B(n13221), .C(n13222), .Y(n4932) );
  INVX1 U11026 ( .A(N3878), .Y(n15503) );
  MUX2X1 U11027 ( .B(n15504), .A(n12626), .S(n13221), .Y(n4931) );
  INVX1 U11028 ( .A(N3874), .Y(n15504) );
  OAI21X1 U11029 ( .A(n15505), .B(n13221), .C(n13222), .Y(n4930) );
  INVX1 U11030 ( .A(N3875), .Y(n15505) );
  MUX2X1 U11031 ( .B(n15506), .A(n12625), .S(n13221), .Y(n4929) );
  INVX1 U11032 ( .A(N3871), .Y(n15506) );
  OAI21X1 U11033 ( .A(n15507), .B(n13221), .C(n13222), .Y(n4928) );
  INVX1 U11034 ( .A(N3872), .Y(n15507) );
  MUX2X1 U11035 ( .B(n15508), .A(n12624), .S(n13221), .Y(n4927) );
  INVX1 U11036 ( .A(N3868), .Y(n15508) );
  OAI21X1 U11037 ( .A(n15509), .B(n13221), .C(n13222), .Y(n4926) );
  NAND2X1 U11038 ( .A(n13221), .B(n12630), .Y(n13222) );
  NOR2X1 U11039 ( .A(n12735), .B(n13220), .Y(n13221) );
  INVX1 U11040 ( .A(N3869), .Y(n15509) );
  MUX2X1 U11041 ( .B(n15510), .A(n12621), .S(n13223), .Y(n4925) );
  INVX1 U11042 ( .A(N3913), .Y(n15510) );
  OAI21X1 U11043 ( .A(n15511), .B(n13223), .C(n13224), .Y(n4924) );
  INVX1 U11044 ( .A(N3914), .Y(n15511) );
  MUX2X1 U11045 ( .B(n15512), .A(n12631), .S(n13223), .Y(n4923) );
  INVX1 U11046 ( .A(N3910), .Y(n15512) );
  OAI21X1 U11047 ( .A(n15513), .B(n13223), .C(n13224), .Y(n4922) );
  INVX1 U11048 ( .A(N3911), .Y(n15513) );
  MUX2X1 U11049 ( .B(n15514), .A(n12629), .S(n13223), .Y(n4921) );
  INVX1 U11050 ( .A(N3907), .Y(n15514) );
  OAI21X1 U11051 ( .A(n15515), .B(n13223), .C(n13224), .Y(n4920) );
  INVX1 U11052 ( .A(N3908), .Y(n15515) );
  MUX2X1 U11053 ( .B(n15516), .A(n12628), .S(n13223), .Y(n4919) );
  INVX1 U11054 ( .A(N3904), .Y(n15516) );
  OAI21X1 U11055 ( .A(n15517), .B(n13223), .C(n13224), .Y(n4918) );
  INVX1 U11056 ( .A(N3905), .Y(n15517) );
  MUX2X1 U11057 ( .B(n15518), .A(n12627), .S(n13223), .Y(n4917) );
  INVX1 U11058 ( .A(N3901), .Y(n15518) );
  OAI21X1 U11059 ( .A(n15519), .B(n13223), .C(n13224), .Y(n4916) );
  INVX1 U11060 ( .A(N3902), .Y(n15519) );
  MUX2X1 U11061 ( .B(n15520), .A(n12626), .S(n13223), .Y(n4915) );
  INVX1 U11062 ( .A(N3898), .Y(n15520) );
  OAI21X1 U11063 ( .A(n15521), .B(n13223), .C(n13224), .Y(n4914) );
  INVX1 U11064 ( .A(N3899), .Y(n15521) );
  MUX2X1 U11065 ( .B(n15522), .A(n12625), .S(n13223), .Y(n4913) );
  INVX1 U11066 ( .A(N3895), .Y(n15522) );
  OAI21X1 U11067 ( .A(n15523), .B(n13223), .C(n13224), .Y(n4912) );
  INVX1 U11068 ( .A(N3896), .Y(n15523) );
  MUX2X1 U11069 ( .B(n15524), .A(n12624), .S(n13223), .Y(n4911) );
  INVX1 U11070 ( .A(N3892), .Y(n15524) );
  OAI21X1 U11071 ( .A(n15525), .B(n13223), .C(n13224), .Y(n4910) );
  NAND2X1 U11072 ( .A(n13223), .B(n12630), .Y(n13224) );
  NOR2X1 U11073 ( .A(n13225), .B(n13220), .Y(n13223) );
  INVX1 U11074 ( .A(N3893), .Y(n15525) );
  MUX2X1 U11075 ( .B(n15526), .A(n12621), .S(n13226), .Y(n4909) );
  INVX1 U11076 ( .A(N3937), .Y(n15526) );
  OAI21X1 U11077 ( .A(n15527), .B(n13226), .C(n13227), .Y(n4908) );
  INVX1 U11078 ( .A(N3938), .Y(n15527) );
  MUX2X1 U11079 ( .B(n15528), .A(n12631), .S(n13226), .Y(n4907) );
  INVX1 U11080 ( .A(N3934), .Y(n15528) );
  OAI21X1 U11081 ( .A(n15529), .B(n13226), .C(n13227), .Y(n4906) );
  INVX1 U11082 ( .A(N3935), .Y(n15529) );
  MUX2X1 U11083 ( .B(n15530), .A(n12629), .S(n13226), .Y(n4905) );
  INVX1 U11084 ( .A(N3931), .Y(n15530) );
  OAI21X1 U11085 ( .A(n15531), .B(n13226), .C(n13227), .Y(n4904) );
  INVX1 U11086 ( .A(N3932), .Y(n15531) );
  MUX2X1 U11087 ( .B(n15532), .A(n12628), .S(n13226), .Y(n4903) );
  INVX1 U11088 ( .A(N3928), .Y(n15532) );
  OAI21X1 U11089 ( .A(n15533), .B(n13226), .C(n13227), .Y(n4902) );
  INVX1 U11090 ( .A(N3929), .Y(n15533) );
  MUX2X1 U11091 ( .B(n15534), .A(n12627), .S(n13226), .Y(n4901) );
  INVX1 U11092 ( .A(N3925), .Y(n15534) );
  OAI21X1 U11093 ( .A(n15535), .B(n13226), .C(n13227), .Y(n4900) );
  INVX1 U11094 ( .A(N3926), .Y(n15535) );
  MUX2X1 U11095 ( .B(n15536), .A(n12626), .S(n13226), .Y(n4899) );
  INVX1 U11096 ( .A(N3922), .Y(n15536) );
  OAI21X1 U11097 ( .A(n15537), .B(n13226), .C(n13227), .Y(n4898) );
  INVX1 U11098 ( .A(N3923), .Y(n15537) );
  MUX2X1 U11099 ( .B(n15538), .A(n12625), .S(n13226), .Y(n4897) );
  INVX1 U11100 ( .A(N3919), .Y(n15538) );
  OAI21X1 U11101 ( .A(n15539), .B(n13226), .C(n13227), .Y(n4896) );
  INVX1 U11102 ( .A(N3920), .Y(n15539) );
  MUX2X1 U11103 ( .B(n15540), .A(n12624), .S(n13226), .Y(n4895) );
  INVX1 U11104 ( .A(N3916), .Y(n15540) );
  OAI21X1 U11105 ( .A(n15541), .B(n13226), .C(n13227), .Y(n4894) );
  NAND2X1 U11106 ( .A(n13226), .B(n12630), .Y(n13227) );
  NOR2X1 U11107 ( .A(n13220), .B(n12678), .Y(n13226) );
  INVX1 U11108 ( .A(N3917), .Y(n15541) );
  MUX2X1 U11109 ( .B(n15542), .A(n12621), .S(n13228), .Y(n4893) );
  INVX1 U11110 ( .A(N3961), .Y(n15542) );
  OAI21X1 U11111 ( .A(n15543), .B(n13228), .C(n13229), .Y(n4892) );
  INVX1 U11112 ( .A(N3962), .Y(n15543) );
  MUX2X1 U11113 ( .B(n15544), .A(n12631), .S(n13228), .Y(n4891) );
  INVX1 U11114 ( .A(N3958), .Y(n15544) );
  OAI21X1 U11115 ( .A(n15545), .B(n13228), .C(n13229), .Y(n4890) );
  INVX1 U11116 ( .A(N3959), .Y(n15545) );
  MUX2X1 U11117 ( .B(n15546), .A(n12629), .S(n13228), .Y(n4889) );
  INVX1 U11118 ( .A(N3955), .Y(n15546) );
  OAI21X1 U11119 ( .A(n15547), .B(n13228), .C(n13229), .Y(n4888) );
  INVX1 U11120 ( .A(N3956), .Y(n15547) );
  MUX2X1 U11121 ( .B(n15548), .A(n12628), .S(n13228), .Y(n4887) );
  INVX1 U11122 ( .A(N3952), .Y(n15548) );
  OAI21X1 U11123 ( .A(n15549), .B(n13228), .C(n13229), .Y(n4886) );
  INVX1 U11124 ( .A(N3953), .Y(n15549) );
  MUX2X1 U11125 ( .B(n15550), .A(n12627), .S(n13228), .Y(n4885) );
  INVX1 U11126 ( .A(N3949), .Y(n15550) );
  OAI21X1 U11127 ( .A(n15551), .B(n13228), .C(n13229), .Y(n4884) );
  INVX1 U11128 ( .A(N3950), .Y(n15551) );
  MUX2X1 U11129 ( .B(n15552), .A(n12626), .S(n13228), .Y(n4883) );
  INVX1 U11130 ( .A(N3946), .Y(n15552) );
  OAI21X1 U11131 ( .A(n15553), .B(n13228), .C(n13229), .Y(n4882) );
  INVX1 U11132 ( .A(N3947), .Y(n15553) );
  MUX2X1 U11133 ( .B(n15554), .A(n12625), .S(n13228), .Y(n4881) );
  INVX1 U11134 ( .A(N3943), .Y(n15554) );
  OAI21X1 U11135 ( .A(n15555), .B(n13228), .C(n13229), .Y(n4880) );
  INVX1 U11136 ( .A(N3944), .Y(n15555) );
  MUX2X1 U11137 ( .B(n15556), .A(n12624), .S(n13228), .Y(n4879) );
  INVX1 U11138 ( .A(N3940), .Y(n15556) );
  OAI21X1 U11139 ( .A(n15557), .B(n13228), .C(n13229), .Y(n4878) );
  NAND2X1 U11140 ( .A(n13228), .B(n12630), .Y(n13229) );
  NOR2X1 U11141 ( .A(n13230), .B(n13220), .Y(n13228) );
  INVX1 U11142 ( .A(N3941), .Y(n15557) );
  MUX2X1 U11143 ( .B(n15558), .A(n12621), .S(n13231), .Y(n4877) );
  INVX1 U11144 ( .A(N3985), .Y(n15558) );
  OAI21X1 U11145 ( .A(n15559), .B(n13231), .C(n13232), .Y(n4876) );
  INVX1 U11146 ( .A(N3986), .Y(n15559) );
  MUX2X1 U11147 ( .B(n15560), .A(n12631), .S(n13231), .Y(n4875) );
  INVX1 U11148 ( .A(N3982), .Y(n15560) );
  OAI21X1 U11149 ( .A(n15561), .B(n13231), .C(n13232), .Y(n4874) );
  INVX1 U11150 ( .A(N3983), .Y(n15561) );
  MUX2X1 U11151 ( .B(n15562), .A(n12629), .S(n13231), .Y(n4873) );
  INVX1 U11152 ( .A(N3979), .Y(n15562) );
  OAI21X1 U11153 ( .A(n15563), .B(n13231), .C(n13232), .Y(n4872) );
  INVX1 U11154 ( .A(N3980), .Y(n15563) );
  MUX2X1 U11155 ( .B(n15564), .A(n12628), .S(n13231), .Y(n4871) );
  INVX1 U11156 ( .A(N3976), .Y(n15564) );
  OAI21X1 U11157 ( .A(n15565), .B(n13231), .C(n13232), .Y(n4870) );
  INVX1 U11158 ( .A(N3977), .Y(n15565) );
  MUX2X1 U11159 ( .B(n15566), .A(n12627), .S(n13231), .Y(n4869) );
  INVX1 U11160 ( .A(N3973), .Y(n15566) );
  OAI21X1 U11161 ( .A(n15567), .B(n13231), .C(n13232), .Y(n4868) );
  INVX1 U11162 ( .A(N3974), .Y(n15567) );
  MUX2X1 U11163 ( .B(n15568), .A(n12626), .S(n13231), .Y(n4867) );
  INVX1 U11164 ( .A(N3970), .Y(n15568) );
  OAI21X1 U11165 ( .A(n15569), .B(n13231), .C(n13232), .Y(n4866) );
  INVX1 U11166 ( .A(N3971), .Y(n15569) );
  MUX2X1 U11167 ( .B(n15570), .A(n12625), .S(n13231), .Y(n4865) );
  INVX1 U11168 ( .A(N3967), .Y(n15570) );
  OAI21X1 U11169 ( .A(n15571), .B(n13231), .C(n13232), .Y(n4864) );
  INVX1 U11170 ( .A(N3968), .Y(n15571) );
  MUX2X1 U11171 ( .B(n15572), .A(n12624), .S(n13231), .Y(n4863) );
  INVX1 U11172 ( .A(N3964), .Y(n15572) );
  OAI21X1 U11173 ( .A(n15573), .B(n13231), .C(n13232), .Y(n4862) );
  NAND2X1 U11174 ( .A(n13231), .B(n12630), .Y(n13232) );
  NOR2X1 U11175 ( .A(n13233), .B(n13220), .Y(n13231) );
  INVX1 U11176 ( .A(N3965), .Y(n15573) );
  MUX2X1 U11177 ( .B(n15574), .A(n12621), .S(n13234), .Y(n4861) );
  INVX1 U11178 ( .A(N4009), .Y(n15574) );
  OAI21X1 U11179 ( .A(n15575), .B(n13234), .C(n13235), .Y(n4860) );
  INVX1 U11180 ( .A(N4010), .Y(n15575) );
  MUX2X1 U11181 ( .B(n15576), .A(n12631), .S(n13234), .Y(n4859) );
  INVX1 U11182 ( .A(N4006), .Y(n15576) );
  OAI21X1 U11183 ( .A(n15577), .B(n13234), .C(n13235), .Y(n4858) );
  INVX1 U11184 ( .A(N4007), .Y(n15577) );
  MUX2X1 U11185 ( .B(n15578), .A(n12629), .S(n13234), .Y(n4857) );
  INVX1 U11186 ( .A(N4003), .Y(n15578) );
  OAI21X1 U11187 ( .A(n15579), .B(n13234), .C(n13235), .Y(n4856) );
  INVX1 U11188 ( .A(N4004), .Y(n15579) );
  MUX2X1 U11189 ( .B(n15580), .A(n12628), .S(n13234), .Y(n4855) );
  INVX1 U11190 ( .A(N4000), .Y(n15580) );
  OAI21X1 U11191 ( .A(n15581), .B(n13234), .C(n13235), .Y(n4854) );
  INVX1 U11192 ( .A(N4001), .Y(n15581) );
  MUX2X1 U11193 ( .B(n15582), .A(n12627), .S(n13234), .Y(n4853) );
  INVX1 U11194 ( .A(N3997), .Y(n15582) );
  OAI21X1 U11195 ( .A(n15583), .B(n13234), .C(n13235), .Y(n4852) );
  INVX1 U11196 ( .A(N3998), .Y(n15583) );
  MUX2X1 U11197 ( .B(n15584), .A(n12626), .S(n13234), .Y(n4851) );
  INVX1 U11198 ( .A(N3994), .Y(n15584) );
  OAI21X1 U11199 ( .A(n15585), .B(n13234), .C(n13235), .Y(n4850) );
  INVX1 U11200 ( .A(N3995), .Y(n15585) );
  MUX2X1 U11201 ( .B(n15586), .A(n12625), .S(n13234), .Y(n4849) );
  INVX1 U11202 ( .A(N3991), .Y(n15586) );
  OAI21X1 U11203 ( .A(n15587), .B(n13234), .C(n13235), .Y(n4848) );
  INVX1 U11204 ( .A(N3992), .Y(n15587) );
  MUX2X1 U11205 ( .B(n15588), .A(n12624), .S(n13234), .Y(n4847) );
  INVX1 U11206 ( .A(N3988), .Y(n15588) );
  OAI21X1 U11207 ( .A(n15589), .B(n13234), .C(n13235), .Y(n4846) );
  NAND2X1 U11208 ( .A(n13234), .B(n12630), .Y(n13235) );
  AND2X1 U11209 ( .A(n12781), .B(n12633), .Y(n13234) );
  INVX1 U11210 ( .A(N3989), .Y(n15589) );
  MUX2X1 U11211 ( .B(n15590), .A(n12621), .S(n13236), .Y(n4845) );
  INVX1 U11212 ( .A(N4177), .Y(n15590) );
  OAI21X1 U11213 ( .A(n15591), .B(n13236), .C(n13237), .Y(n4844) );
  INVX1 U11214 ( .A(N4178), .Y(n15591) );
  MUX2X1 U11215 ( .B(n15592), .A(n12631), .S(n13236), .Y(n4843) );
  INVX1 U11216 ( .A(N4174), .Y(n15592) );
  OAI21X1 U11217 ( .A(n15593), .B(n13236), .C(n13237), .Y(n4842) );
  INVX1 U11218 ( .A(N4175), .Y(n15593) );
  MUX2X1 U11219 ( .B(n15594), .A(n12629), .S(n13236), .Y(n4841) );
  INVX1 U11220 ( .A(N4171), .Y(n15594) );
  OAI21X1 U11221 ( .A(n15595), .B(n13236), .C(n13237), .Y(n4840) );
  INVX1 U11222 ( .A(N4172), .Y(n15595) );
  MUX2X1 U11223 ( .B(n15596), .A(n12628), .S(n13236), .Y(n4839) );
  INVX1 U11224 ( .A(N4168), .Y(n15596) );
  OAI21X1 U11225 ( .A(n15597), .B(n13236), .C(n13237), .Y(n4838) );
  INVX1 U11226 ( .A(N4169), .Y(n15597) );
  MUX2X1 U11227 ( .B(n15598), .A(n12627), .S(n13236), .Y(n4837) );
  INVX1 U11228 ( .A(N4165), .Y(n15598) );
  OAI21X1 U11229 ( .A(n15599), .B(n13236), .C(n13237), .Y(n4836) );
  INVX1 U11230 ( .A(N4166), .Y(n15599) );
  MUX2X1 U11231 ( .B(n15600), .A(n12626), .S(n13236), .Y(n4835) );
  INVX1 U11232 ( .A(N4162), .Y(n15600) );
  OAI21X1 U11233 ( .A(n15601), .B(n13236), .C(n13237), .Y(n4834) );
  INVX1 U11234 ( .A(N4163), .Y(n15601) );
  MUX2X1 U11235 ( .B(n15602), .A(n12625), .S(n13236), .Y(n4833) );
  INVX1 U11236 ( .A(N4159), .Y(n15602) );
  OAI21X1 U11237 ( .A(n15603), .B(n13236), .C(n13237), .Y(n4832) );
  INVX1 U11238 ( .A(N4160), .Y(n15603) );
  MUX2X1 U11239 ( .B(n15604), .A(n12624), .S(n13236), .Y(n4831) );
  INVX1 U11240 ( .A(N4156), .Y(n15604) );
  OAI21X1 U11241 ( .A(n15605), .B(n13236), .C(n13237), .Y(n4830) );
  NAND2X1 U11242 ( .A(n13236), .B(n12630), .Y(n13237) );
  NOR2X1 U11243 ( .A(n13238), .B(n13220), .Y(n13236) );
  INVX1 U11244 ( .A(N4157), .Y(n15605) );
  MUX2X1 U11245 ( .B(n15606), .A(n12621), .S(n13239), .Y(n4829) );
  INVX1 U11246 ( .A(N4201), .Y(n15606) );
  OAI21X1 U11247 ( .A(n15607), .B(n13239), .C(n13240), .Y(n4828) );
  INVX1 U11248 ( .A(N4202), .Y(n15607) );
  MUX2X1 U11249 ( .B(n15608), .A(n12631), .S(n13239), .Y(n4827) );
  INVX1 U11250 ( .A(N4198), .Y(n15608) );
  OAI21X1 U11251 ( .A(n15609), .B(n13239), .C(n13240), .Y(n4826) );
  INVX1 U11252 ( .A(N4199), .Y(n15609) );
  MUX2X1 U11253 ( .B(n15610), .A(n12629), .S(n13239), .Y(n4825) );
  INVX1 U11254 ( .A(N4195), .Y(n15610) );
  OAI21X1 U11255 ( .A(n15611), .B(n13239), .C(n13240), .Y(n4824) );
  INVX1 U11256 ( .A(N4196), .Y(n15611) );
  MUX2X1 U11257 ( .B(n15612), .A(n12628), .S(n13239), .Y(n4823) );
  INVX1 U11258 ( .A(N4192), .Y(n15612) );
  OAI21X1 U11259 ( .A(n15613), .B(n13239), .C(n13240), .Y(n4822) );
  INVX1 U11260 ( .A(N4193), .Y(n15613) );
  MUX2X1 U11261 ( .B(n15614), .A(n12627), .S(n13239), .Y(n4821) );
  INVX1 U11262 ( .A(N4189), .Y(n15614) );
  OAI21X1 U11263 ( .A(n15615), .B(n13239), .C(n13240), .Y(n4820) );
  INVX1 U11264 ( .A(N4190), .Y(n15615) );
  MUX2X1 U11265 ( .B(n15616), .A(n12626), .S(n13239), .Y(n4819) );
  INVX1 U11266 ( .A(N4186), .Y(n15616) );
  OAI21X1 U11267 ( .A(n15617), .B(n13239), .C(n13240), .Y(n4818) );
  INVX1 U11268 ( .A(N4187), .Y(n15617) );
  MUX2X1 U11269 ( .B(n15618), .A(n12625), .S(n13239), .Y(n4817) );
  INVX1 U11270 ( .A(N4183), .Y(n15618) );
  OAI21X1 U11271 ( .A(n15619), .B(n13239), .C(n13240), .Y(n4816) );
  INVX1 U11272 ( .A(N4184), .Y(n15619) );
  MUX2X1 U11273 ( .B(n15620), .A(n12624), .S(n13239), .Y(n4815) );
  INVX1 U11274 ( .A(N4180), .Y(n15620) );
  OAI21X1 U11275 ( .A(n15621), .B(n13239), .C(n13240), .Y(n4814) );
  NAND2X1 U11276 ( .A(n13239), .B(n12630), .Y(n13240) );
  AND2X1 U11277 ( .A(n13241), .B(n12803), .Y(n13239) );
  INVX1 U11278 ( .A(N4181), .Y(n15621) );
  MUX2X1 U11279 ( .B(n12621), .A(n15622), .S(n13242), .Y(n4813) );
  INVX1 U11280 ( .A(N4369), .Y(n15622) );
  OAI21X1 U11281 ( .A(n15623), .B(n13243), .C(n13244), .Y(n4812) );
  INVX1 U11282 ( .A(N4370), .Y(n15623) );
  MUX2X1 U11283 ( .B(n12631), .A(n15624), .S(n13242), .Y(n4811) );
  INVX1 U11284 ( .A(N4366), .Y(n15624) );
  OAI21X1 U11285 ( .A(n15625), .B(n13243), .C(n13244), .Y(n4810) );
  INVX1 U11286 ( .A(N4367), .Y(n15625) );
  MUX2X1 U11287 ( .B(n12629), .A(n15626), .S(n13242), .Y(n4809) );
  INVX1 U11288 ( .A(N4363), .Y(n15626) );
  OAI21X1 U11289 ( .A(n15627), .B(n13243), .C(n13244), .Y(n4808) );
  INVX1 U11290 ( .A(N4364), .Y(n15627) );
  MUX2X1 U11291 ( .B(n12628), .A(n15628), .S(n13242), .Y(n4807) );
  INVX1 U11292 ( .A(N4360), .Y(n15628) );
  OAI21X1 U11293 ( .A(n15629), .B(n13243), .C(n13244), .Y(n4806) );
  INVX1 U11294 ( .A(N4361), .Y(n15629) );
  MUX2X1 U11295 ( .B(n12627), .A(n15630), .S(n13242), .Y(n4805) );
  INVX1 U11296 ( .A(N4357), .Y(n15630) );
  OAI21X1 U11297 ( .A(n15631), .B(n13243), .C(n13244), .Y(n4804) );
  INVX1 U11298 ( .A(N4358), .Y(n15631) );
  MUX2X1 U11299 ( .B(n12626), .A(n15632), .S(n13242), .Y(n4803) );
  INVX1 U11300 ( .A(N4354), .Y(n15632) );
  OAI21X1 U11301 ( .A(n15633), .B(n13243), .C(n13244), .Y(n4802) );
  INVX1 U11302 ( .A(N4355), .Y(n15633) );
  MUX2X1 U11303 ( .B(n12625), .A(n15634), .S(n13242), .Y(n4801) );
  INVX1 U11304 ( .A(N4351), .Y(n15634) );
  OAI21X1 U11305 ( .A(n15635), .B(n13243), .C(n13244), .Y(n4800) );
  INVX1 U11306 ( .A(N4352), .Y(n15635) );
  MUX2X1 U11307 ( .B(n12624), .A(n15636), .S(n13242), .Y(n4799) );
  INVX1 U11308 ( .A(N4348), .Y(n15636) );
  OAI21X1 U11309 ( .A(n15637), .B(n13243), .C(n13244), .Y(n4798) );
  NAND2X1 U11310 ( .A(n13243), .B(n12630), .Y(n13244) );
  INVX1 U11311 ( .A(n13242), .Y(n13243) );
  NAND3X1 U11312 ( .A(n12636), .B(n12816), .C(n12817), .Y(n13242) );
  INVX1 U11313 ( .A(N4349), .Y(n15637) );
  MUX2X1 U11314 ( .B(n15638), .A(n12621), .S(n13245), .Y(n4797) );
  INVX1 U11315 ( .A(N4129), .Y(n15638) );
  OAI21X1 U11316 ( .A(n15639), .B(n13245), .C(n13246), .Y(n4796) );
  INVX1 U11317 ( .A(N4130), .Y(n15639) );
  MUX2X1 U11318 ( .B(n15640), .A(n12631), .S(n13245), .Y(n4795) );
  INVX1 U11319 ( .A(N4126), .Y(n15640) );
  OAI21X1 U11320 ( .A(n15641), .B(n13245), .C(n13246), .Y(n4794) );
  INVX1 U11321 ( .A(N4127), .Y(n15641) );
  MUX2X1 U11322 ( .B(n15642), .A(n12629), .S(n13245), .Y(n4793) );
  INVX1 U11323 ( .A(N4123), .Y(n15642) );
  OAI21X1 U11324 ( .A(n15643), .B(n13245), .C(n13246), .Y(n4792) );
  INVX1 U11325 ( .A(N4124), .Y(n15643) );
  MUX2X1 U11326 ( .B(n15644), .A(n12628), .S(n13245), .Y(n4791) );
  INVX1 U11327 ( .A(N4120), .Y(n15644) );
  OAI21X1 U11328 ( .A(n15645), .B(n13245), .C(n13246), .Y(n4790) );
  INVX1 U11329 ( .A(N4121), .Y(n15645) );
  MUX2X1 U11330 ( .B(n15646), .A(n12627), .S(n13245), .Y(n4789) );
  INVX1 U11331 ( .A(N4117), .Y(n15646) );
  OAI21X1 U11332 ( .A(n15647), .B(n13245), .C(n13246), .Y(n4788) );
  INVX1 U11333 ( .A(N4118), .Y(n15647) );
  MUX2X1 U11334 ( .B(n15648), .A(n12626), .S(n13245), .Y(n4787) );
  INVX1 U11335 ( .A(N4114), .Y(n15648) );
  OAI21X1 U11336 ( .A(n15649), .B(n13245), .C(n13246), .Y(n4786) );
  INVX1 U11337 ( .A(N4115), .Y(n15649) );
  MUX2X1 U11338 ( .B(n15650), .A(n12625), .S(n13245), .Y(n4785) );
  INVX1 U11339 ( .A(N4111), .Y(n15650) );
  OAI21X1 U11340 ( .A(n15651), .B(n13245), .C(n13246), .Y(n4784) );
  INVX1 U11341 ( .A(N4112), .Y(n15651) );
  MUX2X1 U11342 ( .B(n15652), .A(n12624), .S(n13245), .Y(n4783) );
  INVX1 U11343 ( .A(N4108), .Y(n15652) );
  OAI21X1 U11344 ( .A(n15653), .B(n13245), .C(n13246), .Y(n4782) );
  NAND2X1 U11345 ( .A(n13245), .B(n12630), .Y(n13246) );
  AND2X1 U11346 ( .A(n12830), .B(n12633), .Y(n13245) );
  INVX1 U11347 ( .A(n13247), .Y(n12830) );
  INVX1 U11348 ( .A(N4109), .Y(n15653) );
  MUX2X1 U11349 ( .B(n15654), .A(n12621), .S(n13248), .Y(n4781) );
  INVX1 U11350 ( .A(N4153), .Y(n15654) );
  OAI21X1 U11351 ( .A(n15655), .B(n13248), .C(n13249), .Y(n4780) );
  INVX1 U11352 ( .A(N4154), .Y(n15655) );
  MUX2X1 U11353 ( .B(n15656), .A(n12631), .S(n13248), .Y(n4779) );
  INVX1 U11354 ( .A(N4150), .Y(n15656) );
  OAI21X1 U11355 ( .A(n15657), .B(n13248), .C(n13249), .Y(n4778) );
  INVX1 U11356 ( .A(N4151), .Y(n15657) );
  MUX2X1 U11357 ( .B(n15658), .A(n12629), .S(n13248), .Y(n4777) );
  INVX1 U11358 ( .A(N4147), .Y(n15658) );
  OAI21X1 U11359 ( .A(n15659), .B(n13248), .C(n13249), .Y(n4776) );
  INVX1 U11360 ( .A(N4148), .Y(n15659) );
  MUX2X1 U11361 ( .B(n15660), .A(n12628), .S(n13248), .Y(n4775) );
  INVX1 U11362 ( .A(N4144), .Y(n15660) );
  OAI21X1 U11363 ( .A(n15661), .B(n13248), .C(n13249), .Y(n4774) );
  INVX1 U11364 ( .A(N4145), .Y(n15661) );
  MUX2X1 U11365 ( .B(n15662), .A(n12627), .S(n13248), .Y(n4773) );
  INVX1 U11366 ( .A(N4141), .Y(n15662) );
  OAI21X1 U11367 ( .A(n15663), .B(n13248), .C(n13249), .Y(n4772) );
  INVX1 U11368 ( .A(N4142), .Y(n15663) );
  MUX2X1 U11369 ( .B(n15664), .A(n12626), .S(n13248), .Y(n4771) );
  INVX1 U11370 ( .A(N4138), .Y(n15664) );
  OAI21X1 U11371 ( .A(n15665), .B(n13248), .C(n13249), .Y(n4770) );
  INVX1 U11372 ( .A(N4139), .Y(n15665) );
  MUX2X1 U11373 ( .B(n15666), .A(n12625), .S(n13248), .Y(n4769) );
  INVX1 U11374 ( .A(N4135), .Y(n15666) );
  OAI21X1 U11375 ( .A(n15667), .B(n13248), .C(n13249), .Y(n4768) );
  INVX1 U11376 ( .A(N4136), .Y(n15667) );
  MUX2X1 U11377 ( .B(n15668), .A(n12624), .S(n13248), .Y(n4767) );
  INVX1 U11378 ( .A(N4132), .Y(n15668) );
  OAI21X1 U11379 ( .A(n15669), .B(n13248), .C(n13249), .Y(n4766) );
  NAND2X1 U11380 ( .A(n13248), .B(n12630), .Y(n13249) );
  AND2X1 U11381 ( .A(n12633), .B(n13250), .Y(n13248) );
  INVX1 U11382 ( .A(N4133), .Y(n15669) );
  MUX2X1 U11383 ( .B(n15670), .A(n12621), .S(n13251), .Y(n4765) );
  INVX1 U11384 ( .A(N4321), .Y(n15670) );
  OAI21X1 U11385 ( .A(n15671), .B(n13251), .C(n13252), .Y(n4764) );
  INVX1 U11386 ( .A(N4322), .Y(n15671) );
  MUX2X1 U11387 ( .B(n15672), .A(n12631), .S(n13251), .Y(n4763) );
  INVX1 U11388 ( .A(N4318), .Y(n15672) );
  OAI21X1 U11389 ( .A(n15673), .B(n13251), .C(n13252), .Y(n4762) );
  INVX1 U11390 ( .A(N4319), .Y(n15673) );
  MUX2X1 U11391 ( .B(n15674), .A(n12629), .S(n13251), .Y(n4761) );
  INVX1 U11392 ( .A(N4315), .Y(n15674) );
  OAI21X1 U11393 ( .A(n15675), .B(n13251), .C(n13252), .Y(n4760) );
  INVX1 U11394 ( .A(N4316), .Y(n15675) );
  MUX2X1 U11395 ( .B(n15676), .A(n12628), .S(n13251), .Y(n4759) );
  INVX1 U11396 ( .A(N4312), .Y(n15676) );
  OAI21X1 U11397 ( .A(n15677), .B(n13251), .C(n13252), .Y(n4758) );
  INVX1 U11398 ( .A(N4313), .Y(n15677) );
  MUX2X1 U11399 ( .B(n15678), .A(n12627), .S(n13251), .Y(n4757) );
  INVX1 U11400 ( .A(N4309), .Y(n15678) );
  OAI21X1 U11401 ( .A(n15679), .B(n13251), .C(n13252), .Y(n4756) );
  INVX1 U11402 ( .A(N4310), .Y(n15679) );
  MUX2X1 U11403 ( .B(n15680), .A(n12626), .S(n13251), .Y(n4755) );
  INVX1 U11404 ( .A(N4306), .Y(n15680) );
  OAI21X1 U11405 ( .A(n15681), .B(n13251), .C(n13252), .Y(n4754) );
  INVX1 U11406 ( .A(N4307), .Y(n15681) );
  MUX2X1 U11407 ( .B(n15682), .A(n12625), .S(n13251), .Y(n4753) );
  INVX1 U11408 ( .A(N4303), .Y(n15682) );
  OAI21X1 U11409 ( .A(n15683), .B(n13251), .C(n13252), .Y(n4752) );
  INVX1 U11410 ( .A(N4304), .Y(n15683) );
  MUX2X1 U11411 ( .B(n15684), .A(n12624), .S(n13251), .Y(n4751) );
  INVX1 U11412 ( .A(N4300), .Y(n15684) );
  OAI21X1 U11413 ( .A(n15685), .B(n13251), .C(n13252), .Y(n4750) );
  NAND2X1 U11414 ( .A(n13251), .B(n12630), .Y(n13252) );
  AND2X1 U11415 ( .A(n13241), .B(n12841), .Y(n13251) );
  INVX1 U11416 ( .A(n13253), .Y(n12841) );
  INVX1 U11417 ( .A(N4301), .Y(n15685) );
  MUX2X1 U11418 ( .B(n15686), .A(n12621), .S(n13254), .Y(n4749) );
  INVX1 U11419 ( .A(N4345), .Y(n15686) );
  OAI21X1 U11420 ( .A(n15687), .B(n13254), .C(n13255), .Y(n4748) );
  INVX1 U11421 ( .A(N4346), .Y(n15687) );
  MUX2X1 U11422 ( .B(n15688), .A(n12631), .S(n13254), .Y(n4747) );
  INVX1 U11423 ( .A(N4342), .Y(n15688) );
  OAI21X1 U11424 ( .A(n15689), .B(n13254), .C(n13255), .Y(n4746) );
  INVX1 U11425 ( .A(N4343), .Y(n15689) );
  MUX2X1 U11426 ( .B(n15690), .A(n12629), .S(n13254), .Y(n4745) );
  INVX1 U11427 ( .A(N4339), .Y(n15690) );
  OAI21X1 U11428 ( .A(n15691), .B(n13254), .C(n13255), .Y(n4744) );
  INVX1 U11429 ( .A(N4340), .Y(n15691) );
  MUX2X1 U11430 ( .B(n15692), .A(n12628), .S(n13254), .Y(n4743) );
  INVX1 U11431 ( .A(N4336), .Y(n15692) );
  OAI21X1 U11432 ( .A(n15693), .B(n13254), .C(n13255), .Y(n4742) );
  INVX1 U11433 ( .A(N4337), .Y(n15693) );
  MUX2X1 U11434 ( .B(n15694), .A(n12627), .S(n13254), .Y(n4741) );
  INVX1 U11435 ( .A(N4333), .Y(n15694) );
  OAI21X1 U11436 ( .A(n15695), .B(n13254), .C(n13255), .Y(n4740) );
  INVX1 U11437 ( .A(N4334), .Y(n15695) );
  MUX2X1 U11438 ( .B(n15696), .A(n12626), .S(n13254), .Y(n4739) );
  INVX1 U11439 ( .A(N4330), .Y(n15696) );
  OAI21X1 U11440 ( .A(n15697), .B(n13254), .C(n13255), .Y(n4738) );
  INVX1 U11441 ( .A(N4331), .Y(n15697) );
  MUX2X1 U11442 ( .B(n15698), .A(n12625), .S(n13254), .Y(n4737) );
  INVX1 U11443 ( .A(N4327), .Y(n15698) );
  OAI21X1 U11444 ( .A(n15699), .B(n13254), .C(n13255), .Y(n4736) );
  INVX1 U11445 ( .A(N4328), .Y(n15699) );
  MUX2X1 U11446 ( .B(n15700), .A(n12624), .S(n13254), .Y(n4735) );
  INVX1 U11447 ( .A(N4324), .Y(n15700) );
  OAI21X1 U11448 ( .A(n15701), .B(n13254), .C(n13255), .Y(n4734) );
  NAND2X1 U11449 ( .A(n13254), .B(n12630), .Y(n13255) );
  AND2X1 U11450 ( .A(n13241), .B(n12851), .Y(n13254) );
  INVX1 U11451 ( .A(n13256), .Y(n12851) );
  INVX1 U11452 ( .A(N4325), .Y(n15701) );
  MUX2X1 U11453 ( .B(n15702), .A(n12621), .S(n13257), .Y(n4733) );
  INVX1 U11454 ( .A(N4105), .Y(n15702) );
  OAI21X1 U11455 ( .A(n15703), .B(n13257), .C(n13258), .Y(n4732) );
  INVX1 U11456 ( .A(N4106), .Y(n15703) );
  MUX2X1 U11457 ( .B(n15704), .A(n12631), .S(n13257), .Y(n4731) );
  INVX1 U11458 ( .A(N4102), .Y(n15704) );
  OAI21X1 U11459 ( .A(n15705), .B(n13257), .C(n13258), .Y(n4730) );
  INVX1 U11460 ( .A(N4103), .Y(n15705) );
  MUX2X1 U11461 ( .B(n15706), .A(n12629), .S(n13257), .Y(n4729) );
  INVX1 U11462 ( .A(N4099), .Y(n15706) );
  OAI21X1 U11463 ( .A(n15707), .B(n13257), .C(n13258), .Y(n4728) );
  INVX1 U11464 ( .A(N4100), .Y(n15707) );
  MUX2X1 U11465 ( .B(n15708), .A(n12628), .S(n13257), .Y(n4727) );
  INVX1 U11466 ( .A(N4096), .Y(n15708) );
  OAI21X1 U11467 ( .A(n15709), .B(n13257), .C(n13258), .Y(n4726) );
  INVX1 U11468 ( .A(N4097), .Y(n15709) );
  MUX2X1 U11469 ( .B(n15710), .A(n12627), .S(n13257), .Y(n4725) );
  INVX1 U11470 ( .A(N4093), .Y(n15710) );
  OAI21X1 U11471 ( .A(n15711), .B(n13257), .C(n13258), .Y(n4724) );
  INVX1 U11472 ( .A(N4094), .Y(n15711) );
  MUX2X1 U11473 ( .B(n15712), .A(n12626), .S(n13257), .Y(n4723) );
  INVX1 U11474 ( .A(N4090), .Y(n15712) );
  OAI21X1 U11475 ( .A(n15713), .B(n13257), .C(n13258), .Y(n4722) );
  INVX1 U11476 ( .A(N4091), .Y(n15713) );
  MUX2X1 U11477 ( .B(n15714), .A(n12625), .S(n13257), .Y(n4721) );
  INVX1 U11478 ( .A(N4087), .Y(n15714) );
  OAI21X1 U11479 ( .A(n15715), .B(n13257), .C(n13258), .Y(n4720) );
  INVX1 U11480 ( .A(N4088), .Y(n15715) );
  MUX2X1 U11481 ( .B(n15716), .A(n12624), .S(n13257), .Y(n4719) );
  INVX1 U11482 ( .A(N4084), .Y(n15716) );
  OAI21X1 U11483 ( .A(n15717), .B(n13257), .C(n13258), .Y(n4718) );
  NAND2X1 U11484 ( .A(n13257), .B(n12630), .Y(n13258) );
  AND2X1 U11485 ( .A(n12633), .B(n13259), .Y(n13257) );
  INVX1 U11486 ( .A(N4085), .Y(n15717) );
  MUX2X1 U11487 ( .B(n15718), .A(n12621), .S(n13260), .Y(n4717) );
  INVX1 U11488 ( .A(N4273), .Y(n15718) );
  OAI21X1 U11489 ( .A(n15719), .B(n13260), .C(n13261), .Y(n4716) );
  INVX1 U11490 ( .A(N4274), .Y(n15719) );
  MUX2X1 U11491 ( .B(n15720), .A(n12631), .S(n13260), .Y(n4715) );
  INVX1 U11492 ( .A(N4270), .Y(n15720) );
  OAI21X1 U11493 ( .A(n15721), .B(n13260), .C(n13261), .Y(n4714) );
  INVX1 U11494 ( .A(N4271), .Y(n15721) );
  MUX2X1 U11495 ( .B(n15722), .A(n12629), .S(n13260), .Y(n4713) );
  INVX1 U11496 ( .A(N4267), .Y(n15722) );
  OAI21X1 U11497 ( .A(n15723), .B(n13260), .C(n13261), .Y(n4712) );
  INVX1 U11498 ( .A(N4268), .Y(n15723) );
  MUX2X1 U11499 ( .B(n15724), .A(n12628), .S(n13260), .Y(n4711) );
  INVX1 U11500 ( .A(N4264), .Y(n15724) );
  OAI21X1 U11501 ( .A(n15725), .B(n13260), .C(n13261), .Y(n4710) );
  INVX1 U11502 ( .A(N4265), .Y(n15725) );
  MUX2X1 U11503 ( .B(n15726), .A(n12627), .S(n13260), .Y(n4709) );
  INVX1 U11504 ( .A(N4261), .Y(n15726) );
  OAI21X1 U11505 ( .A(n15727), .B(n13260), .C(n13261), .Y(n4708) );
  INVX1 U11506 ( .A(N4262), .Y(n15727) );
  MUX2X1 U11507 ( .B(n15728), .A(n12626), .S(n13260), .Y(n4707) );
  INVX1 U11508 ( .A(N4258), .Y(n15728) );
  OAI21X1 U11509 ( .A(n15729), .B(n13260), .C(n13261), .Y(n4706) );
  INVX1 U11510 ( .A(N4259), .Y(n15729) );
  MUX2X1 U11511 ( .B(n15730), .A(n12625), .S(n13260), .Y(n4705) );
  INVX1 U11512 ( .A(N4255), .Y(n15730) );
  OAI21X1 U11513 ( .A(n15731), .B(n13260), .C(n13261), .Y(n4704) );
  INVX1 U11514 ( .A(N4256), .Y(n15731) );
  MUX2X1 U11515 ( .B(n15732), .A(n12624), .S(n13260), .Y(n4703) );
  INVX1 U11516 ( .A(N4252), .Y(n15732) );
  OAI21X1 U11517 ( .A(n15733), .B(n13260), .C(n13261), .Y(n4702) );
  NAND2X1 U11518 ( .A(n13260), .B(n12630), .Y(n13261) );
  AND2X1 U11519 ( .A(n13241), .B(n12870), .Y(n13260) );
  INVX1 U11520 ( .A(N4253), .Y(n15733) );
  MUX2X1 U11521 ( .B(n15734), .A(n12621), .S(n13262), .Y(n4701) );
  INVX1 U11522 ( .A(N4297), .Y(n15734) );
  OAI21X1 U11523 ( .A(n15735), .B(n13262), .C(n13263), .Y(n4700) );
  INVX1 U11524 ( .A(N4298), .Y(n15735) );
  MUX2X1 U11525 ( .B(n15736), .A(n12631), .S(n13262), .Y(n4699) );
  INVX1 U11526 ( .A(N4294), .Y(n15736) );
  OAI21X1 U11527 ( .A(n15737), .B(n13262), .C(n13263), .Y(n4698) );
  INVX1 U11528 ( .A(N4295), .Y(n15737) );
  MUX2X1 U11529 ( .B(n15738), .A(n12629), .S(n13262), .Y(n4697) );
  INVX1 U11530 ( .A(N4291), .Y(n15738) );
  OAI21X1 U11531 ( .A(n15739), .B(n13262), .C(n13263), .Y(n4696) );
  INVX1 U11532 ( .A(N4292), .Y(n15739) );
  MUX2X1 U11533 ( .B(n15740), .A(n12628), .S(n13262), .Y(n4695) );
  INVX1 U11534 ( .A(N4288), .Y(n15740) );
  OAI21X1 U11535 ( .A(n15741), .B(n13262), .C(n13263), .Y(n4694) );
  INVX1 U11536 ( .A(N4289), .Y(n15741) );
  MUX2X1 U11537 ( .B(n15742), .A(n12627), .S(n13262), .Y(n4693) );
  INVX1 U11538 ( .A(N4285), .Y(n15742) );
  OAI21X1 U11539 ( .A(n15743), .B(n13262), .C(n13263), .Y(n4692) );
  INVX1 U11540 ( .A(N4286), .Y(n15743) );
  MUX2X1 U11541 ( .B(n15744), .A(n12626), .S(n13262), .Y(n4691) );
  INVX1 U11542 ( .A(N4282), .Y(n15744) );
  OAI21X1 U11543 ( .A(n15745), .B(n13262), .C(n13263), .Y(n4690) );
  INVX1 U11544 ( .A(N4283), .Y(n15745) );
  MUX2X1 U11545 ( .B(n15746), .A(n12625), .S(n13262), .Y(n4689) );
  INVX1 U11546 ( .A(N4279), .Y(n15746) );
  OAI21X1 U11547 ( .A(n15747), .B(n13262), .C(n13263), .Y(n4688) );
  INVX1 U11548 ( .A(N4280), .Y(n15747) );
  MUX2X1 U11549 ( .B(n15748), .A(n12624), .S(n13262), .Y(n4687) );
  INVX1 U11550 ( .A(N4276), .Y(n15748) );
  OAI21X1 U11551 ( .A(n15749), .B(n13262), .C(n13263), .Y(n4686) );
  NAND2X1 U11552 ( .A(n13262), .B(n12630), .Y(n13263) );
  AND2X1 U11553 ( .A(n13241), .B(n12880), .Y(n13262) );
  INVX1 U11554 ( .A(N4277), .Y(n15749) );
  MUX2X1 U11555 ( .B(n15750), .A(n12621), .S(n13264), .Y(n4685) );
  INVX1 U11556 ( .A(N4033), .Y(n15750) );
  OAI21X1 U11557 ( .A(n15751), .B(n13264), .C(n13265), .Y(n4684) );
  INVX1 U11558 ( .A(N4034), .Y(n15751) );
  MUX2X1 U11559 ( .B(n15752), .A(n12631), .S(n13264), .Y(n4683) );
  INVX1 U11560 ( .A(N4030), .Y(n15752) );
  OAI21X1 U11561 ( .A(n15753), .B(n13264), .C(n13265), .Y(n4682) );
  INVX1 U11562 ( .A(N4031), .Y(n15753) );
  MUX2X1 U11563 ( .B(n15754), .A(n12629), .S(n13264), .Y(n4681) );
  INVX1 U11564 ( .A(N4027), .Y(n15754) );
  OAI21X1 U11565 ( .A(n15755), .B(n13264), .C(n13265), .Y(n4680) );
  INVX1 U11566 ( .A(N4028), .Y(n15755) );
  MUX2X1 U11567 ( .B(n15756), .A(n12628), .S(n13264), .Y(n4679) );
  INVX1 U11568 ( .A(N4024), .Y(n15756) );
  OAI21X1 U11569 ( .A(n15757), .B(n13264), .C(n13265), .Y(n4678) );
  INVX1 U11570 ( .A(N4025), .Y(n15757) );
  MUX2X1 U11571 ( .B(n15758), .A(n12627), .S(n13264), .Y(n4677) );
  INVX1 U11572 ( .A(N4021), .Y(n15758) );
  OAI21X1 U11573 ( .A(n15759), .B(n13264), .C(n13265), .Y(n4676) );
  INVX1 U11574 ( .A(N4022), .Y(n15759) );
  MUX2X1 U11575 ( .B(n15760), .A(n12626), .S(n13264), .Y(n4675) );
  INVX1 U11576 ( .A(N4018), .Y(n15760) );
  OAI21X1 U11577 ( .A(n15761), .B(n13264), .C(n13265), .Y(n4674) );
  INVX1 U11578 ( .A(N4019), .Y(n15761) );
  MUX2X1 U11579 ( .B(n15762), .A(n12625), .S(n13264), .Y(n4673) );
  INVX1 U11580 ( .A(N4015), .Y(n15762) );
  OAI21X1 U11581 ( .A(n15763), .B(n13264), .C(n13265), .Y(n4672) );
  INVX1 U11582 ( .A(N4016), .Y(n15763) );
  MUX2X1 U11583 ( .B(n15764), .A(n12624), .S(n13264), .Y(n4671) );
  INVX1 U11584 ( .A(N4012), .Y(n15764) );
  OAI21X1 U11585 ( .A(n15765), .B(n13264), .C(n13265), .Y(n4670) );
  NAND2X1 U11586 ( .A(n13264), .B(n12630), .Y(n13265) );
  AND2X1 U11587 ( .A(n12890), .B(n12633), .Y(n13264) );
  INVX1 U11588 ( .A(N4013), .Y(n15765) );
  MUX2X1 U11589 ( .B(n15766), .A(n12621), .S(n13266), .Y(n4669) );
  INVX1 U11590 ( .A(N4057), .Y(n15766) );
  OAI21X1 U11591 ( .A(n15767), .B(n13266), .C(n13267), .Y(n4668) );
  INVX1 U11592 ( .A(N4058), .Y(n15767) );
  MUX2X1 U11593 ( .B(n15768), .A(n12631), .S(n13266), .Y(n4667) );
  INVX1 U11594 ( .A(N4054), .Y(n15768) );
  OAI21X1 U11595 ( .A(n15769), .B(n13266), .C(n13267), .Y(n4666) );
  INVX1 U11596 ( .A(N4055), .Y(n15769) );
  MUX2X1 U11597 ( .B(n15770), .A(n12629), .S(n13266), .Y(n4665) );
  INVX1 U11598 ( .A(N4051), .Y(n15770) );
  OAI21X1 U11599 ( .A(n15771), .B(n13266), .C(n13267), .Y(n4664) );
  INVX1 U11600 ( .A(N4052), .Y(n15771) );
  MUX2X1 U11601 ( .B(n15772), .A(n12628), .S(n13266), .Y(n4663) );
  INVX1 U11602 ( .A(N4048), .Y(n15772) );
  OAI21X1 U11603 ( .A(n15773), .B(n13266), .C(n13267), .Y(n4662) );
  INVX1 U11604 ( .A(N4049), .Y(n15773) );
  MUX2X1 U11605 ( .B(n15774), .A(n12627), .S(n13266), .Y(n4661) );
  INVX1 U11606 ( .A(N4045), .Y(n15774) );
  OAI21X1 U11607 ( .A(n15775), .B(n13266), .C(n13267), .Y(n4660) );
  INVX1 U11608 ( .A(N4046), .Y(n15775) );
  MUX2X1 U11609 ( .B(n15776), .A(n12626), .S(n13266), .Y(n4659) );
  INVX1 U11610 ( .A(N4042), .Y(n15776) );
  OAI21X1 U11611 ( .A(n15777), .B(n13266), .C(n13267), .Y(n4658) );
  INVX1 U11612 ( .A(N4043), .Y(n15777) );
  MUX2X1 U11613 ( .B(n15778), .A(n12625), .S(n13266), .Y(n4657) );
  INVX1 U11614 ( .A(N4039), .Y(n15778) );
  OAI21X1 U11615 ( .A(n15779), .B(n13266), .C(n13267), .Y(n4656) );
  INVX1 U11616 ( .A(N4040), .Y(n15779) );
  MUX2X1 U11617 ( .B(n15780), .A(n12624), .S(n13266), .Y(n4655) );
  INVX1 U11618 ( .A(N4036), .Y(n15780) );
  OAI21X1 U11619 ( .A(n15781), .B(n13266), .C(n13267), .Y(n4654) );
  NAND2X1 U11620 ( .A(n13266), .B(n12630), .Y(n13267) );
  AND2X1 U11621 ( .A(n12900), .B(n12633), .Y(n13266) );
  NOR2X1 U11622 ( .A(n13220), .B(N981), .Y(n12633) );
  INVX1 U11623 ( .A(n13268), .Y(n12900) );
  INVX1 U11624 ( .A(N4037), .Y(n15781) );
  MUX2X1 U11625 ( .B(n15782), .A(n12621), .S(n13269), .Y(n4653) );
  INVX1 U11626 ( .A(N4225), .Y(n15782) );
  OAI21X1 U11627 ( .A(n15783), .B(n13269), .C(n13270), .Y(n4652) );
  INVX1 U11628 ( .A(N4226), .Y(n15783) );
  MUX2X1 U11629 ( .B(n15784), .A(n12631), .S(n13269), .Y(n4651) );
  INVX1 U11630 ( .A(N4222), .Y(n15784) );
  OAI21X1 U11631 ( .A(n15785), .B(n13269), .C(n13270), .Y(n4650) );
  INVX1 U11632 ( .A(N4223), .Y(n15785) );
  MUX2X1 U11633 ( .B(n15786), .A(n12629), .S(n13269), .Y(n4649) );
  INVX1 U11634 ( .A(N4219), .Y(n15786) );
  OAI21X1 U11635 ( .A(n15787), .B(n13269), .C(n13270), .Y(n4648) );
  INVX1 U11636 ( .A(N4220), .Y(n15787) );
  MUX2X1 U11637 ( .B(n15788), .A(n12628), .S(n13269), .Y(n4647) );
  INVX1 U11638 ( .A(N4216), .Y(n15788) );
  OAI21X1 U11639 ( .A(n15789), .B(n13269), .C(n13270), .Y(n4646) );
  INVX1 U11640 ( .A(N4217), .Y(n15789) );
  MUX2X1 U11641 ( .B(n15790), .A(n12627), .S(n13269), .Y(n4645) );
  INVX1 U11642 ( .A(N4213), .Y(n15790) );
  OAI21X1 U11643 ( .A(n15791), .B(n13269), .C(n13270), .Y(n4644) );
  INVX1 U11644 ( .A(N4214), .Y(n15791) );
  MUX2X1 U11645 ( .B(n15792), .A(n12626), .S(n13269), .Y(n4643) );
  INVX1 U11646 ( .A(N4210), .Y(n15792) );
  OAI21X1 U11647 ( .A(n15793), .B(n13269), .C(n13270), .Y(n4642) );
  INVX1 U11648 ( .A(N4211), .Y(n15793) );
  MUX2X1 U11649 ( .B(n15794), .A(n12625), .S(n13269), .Y(n4641) );
  INVX1 U11650 ( .A(N4207), .Y(n15794) );
  OAI21X1 U11651 ( .A(n15795), .B(n13269), .C(n13270), .Y(n4640) );
  INVX1 U11652 ( .A(N4208), .Y(n15795) );
  MUX2X1 U11653 ( .B(n15796), .A(n12624), .S(n13269), .Y(n4639) );
  INVX1 U11654 ( .A(N4204), .Y(n15796) );
  OAI21X1 U11655 ( .A(n15797), .B(n13269), .C(n13270), .Y(n4638) );
  NAND2X1 U11656 ( .A(n13269), .B(n12630), .Y(n13270) );
  AND2X1 U11657 ( .A(n13241), .B(n13175), .Y(n13269) );
  INVX1 U11658 ( .A(n13271), .Y(n13175) );
  INVX1 U11659 ( .A(N4205), .Y(n15797) );
  MUX2X1 U11660 ( .B(n15798), .A(n12621), .S(n13272), .Y(n4637) );
  INVX1 U11661 ( .A(N4249), .Y(n15798) );
  OAI21X1 U11662 ( .A(n15799), .B(n13272), .C(n13273), .Y(n4636) );
  INVX1 U11663 ( .A(N4250), .Y(n15799) );
  MUX2X1 U11664 ( .B(n15800), .A(n12631), .S(n13272), .Y(n4635) );
  INVX1 U11665 ( .A(N4246), .Y(n15800) );
  OAI21X1 U11666 ( .A(n15801), .B(n13272), .C(n13273), .Y(n4634) );
  INVX1 U11667 ( .A(N4247), .Y(n15801) );
  MUX2X1 U11668 ( .B(n15802), .A(n12629), .S(n13272), .Y(n4633) );
  INVX1 U11669 ( .A(N4243), .Y(n15802) );
  OAI21X1 U11670 ( .A(n15803), .B(n13272), .C(n13273), .Y(n4632) );
  INVX1 U11671 ( .A(N4244), .Y(n15803) );
  MUX2X1 U11672 ( .B(n15804), .A(n12628), .S(n13272), .Y(n4631) );
  INVX1 U11673 ( .A(N4240), .Y(n15804) );
  OAI21X1 U11674 ( .A(n15805), .B(n13272), .C(n13273), .Y(n4630) );
  INVX1 U11675 ( .A(N4241), .Y(n15805) );
  MUX2X1 U11676 ( .B(n15806), .A(n12627), .S(n13272), .Y(n4629) );
  INVX1 U11677 ( .A(N4237), .Y(n15806) );
  OAI21X1 U11678 ( .A(n15807), .B(n13272), .C(n13273), .Y(n4628) );
  INVX1 U11679 ( .A(N4238), .Y(n15807) );
  MUX2X1 U11680 ( .B(n15808), .A(n12626), .S(n13272), .Y(n4627) );
  INVX1 U11681 ( .A(N4234), .Y(n15808) );
  OAI21X1 U11682 ( .A(n15809), .B(n13272), .C(n13273), .Y(n4626) );
  INVX1 U11683 ( .A(N4235), .Y(n15809) );
  MUX2X1 U11684 ( .B(n15810), .A(n12625), .S(n13272), .Y(n4625) );
  INVX1 U11685 ( .A(N4231), .Y(n15810) );
  OAI21X1 U11686 ( .A(n15811), .B(n13272), .C(n13273), .Y(n4624) );
  INVX1 U11687 ( .A(N4232), .Y(n15811) );
  MUX2X1 U11688 ( .B(n15812), .A(n12624), .S(n13272), .Y(n4623) );
  INVX1 U11689 ( .A(N4228), .Y(n15812) );
  OAI21X1 U11690 ( .A(n15813), .B(n13272), .C(n13273), .Y(n4622) );
  NAND2X1 U11691 ( .A(n13272), .B(n12630), .Y(n13273) );
  AND2X1 U11692 ( .A(n13241), .B(n13185), .Y(n13272) );
  NOR2X1 U11693 ( .A(n13220), .B(N980), .Y(n13241) );
  INVX1 U11694 ( .A(N4229), .Y(n15813) );
  OAI21X1 U11695 ( .A(n15814), .B(n13274), .C(n13275), .Y(n4621) );
  INVX1 U11696 ( .A(N3821), .Y(n15814) );
  MUX2X1 U11697 ( .B(n15815), .A(n12624), .S(n13274), .Y(n4620) );
  INVX1 U11698 ( .A(N3820), .Y(n15815) );
  OAI21X1 U11699 ( .A(n15816), .B(n13274), .C(n13275), .Y(n4619) );
  INVX1 U11700 ( .A(N3824), .Y(n15816) );
  MUX2X1 U11701 ( .B(n15817), .A(n12625), .S(n13274), .Y(n4618) );
  INVX1 U11702 ( .A(N3823), .Y(n15817) );
  OAI21X1 U11703 ( .A(n15818), .B(n13274), .C(n13275), .Y(n4617) );
  INVX1 U11704 ( .A(N3827), .Y(n15818) );
  MUX2X1 U11705 ( .B(n15819), .A(n12626), .S(n13274), .Y(n4616) );
  INVX1 U11706 ( .A(N3826), .Y(n15819) );
  OAI21X1 U11707 ( .A(n15820), .B(n13274), .C(n13275), .Y(n4615) );
  INVX1 U11708 ( .A(N3830), .Y(n15820) );
  MUX2X1 U11709 ( .B(n15821), .A(n12627), .S(n13274), .Y(n4614) );
  INVX1 U11710 ( .A(N3829), .Y(n15821) );
  OAI21X1 U11711 ( .A(n15822), .B(n13274), .C(n13275), .Y(n4613) );
  INVX1 U11712 ( .A(N3833), .Y(n15822) );
  MUX2X1 U11713 ( .B(n15823), .A(n12628), .S(n13274), .Y(n4612) );
  INVX1 U11714 ( .A(N3832), .Y(n15823) );
  OAI21X1 U11715 ( .A(n15824), .B(n13274), .C(n13275), .Y(n4611) );
  INVX1 U11716 ( .A(N3836), .Y(n15824) );
  MUX2X1 U11717 ( .B(n15825), .A(n12629), .S(n13274), .Y(n4610) );
  INVX1 U11718 ( .A(N3835), .Y(n15825) );
  OAI21X1 U11719 ( .A(n15826), .B(n13274), .C(n13275), .Y(n4609) );
  INVX1 U11720 ( .A(N3839), .Y(n15826) );
  MUX2X1 U11721 ( .B(n15827), .A(n12631), .S(n13274), .Y(n4608) );
  INVX1 U11722 ( .A(N3838), .Y(n15827) );
  OAI21X1 U11723 ( .A(n15828), .B(n13274), .C(n13275), .Y(n4607) );
  NAND2X1 U11724 ( .A(n13274), .B(n12630), .Y(n13275) );
  INVX1 U11725 ( .A(N3842), .Y(n15828) );
  MUX2X1 U11726 ( .B(n15829), .A(n12621), .S(n13274), .Y(n4606) );
  NOR2X1 U11727 ( .A(n13276), .B(n13220), .Y(n13274) );
  INVX1 U11728 ( .A(N3841), .Y(n15829) );
  OAI21X1 U11729 ( .A(n15830), .B(n13277), .C(n13278), .Y(n4605) );
  INVX1 U11730 ( .A(N3797), .Y(n15830) );
  MUX2X1 U11731 ( .B(n15831), .A(n12624), .S(n13277), .Y(n4604) );
  NAND2X1 U11732 ( .A(n13279), .B(InData[7]), .Y(n12624) );
  INVX1 U11733 ( .A(N3796), .Y(n15831) );
  OAI21X1 U11734 ( .A(n15832), .B(n13277), .C(n13278), .Y(n4603) );
  INVX1 U11735 ( .A(N3800), .Y(n15832) );
  MUX2X1 U11736 ( .B(n15833), .A(n12625), .S(n13277), .Y(n4602) );
  NAND2X1 U11737 ( .A(n13279), .B(InData[6]), .Y(n12625) );
  INVX1 U11738 ( .A(N3799), .Y(n15833) );
  OAI21X1 U11739 ( .A(n15834), .B(n13277), .C(n13278), .Y(n4601) );
  INVX1 U11740 ( .A(N3803), .Y(n15834) );
  MUX2X1 U11741 ( .B(n15835), .A(n12626), .S(n13277), .Y(n4600) );
  NAND2X1 U11742 ( .A(n13279), .B(InData[5]), .Y(n12626) );
  INVX1 U11743 ( .A(N3802), .Y(n15835) );
  OAI21X1 U11744 ( .A(n15836), .B(n13277), .C(n13278), .Y(n4599) );
  INVX1 U11745 ( .A(N3806), .Y(n15836) );
  MUX2X1 U11746 ( .B(n15837), .A(n12627), .S(n13277), .Y(n4598) );
  NAND2X1 U11747 ( .A(n13279), .B(InData[4]), .Y(n12627) );
  INVX1 U11748 ( .A(N3805), .Y(n15837) );
  OAI21X1 U11749 ( .A(n15838), .B(n13277), .C(n13278), .Y(n4597) );
  INVX1 U11750 ( .A(N3809), .Y(n15838) );
  MUX2X1 U11751 ( .B(n15839), .A(n12628), .S(n13277), .Y(n4596) );
  NAND2X1 U11752 ( .A(n13279), .B(InData[3]), .Y(n12628) );
  INVX1 U11753 ( .A(N3808), .Y(n15839) );
  OAI21X1 U11754 ( .A(n15840), .B(n13277), .C(n13278), .Y(n4595) );
  INVX1 U11755 ( .A(N3812), .Y(n15840) );
  MUX2X1 U11756 ( .B(n15841), .A(n12629), .S(n13277), .Y(n4594) );
  NAND2X1 U11757 ( .A(n13279), .B(InData[2]), .Y(n12629) );
  INVX1 U11758 ( .A(N3811), .Y(n15841) );
  OAI21X1 U11759 ( .A(n15842), .B(n13277), .C(n13278), .Y(n4593) );
  INVX1 U11760 ( .A(N3815), .Y(n15842) );
  MUX2X1 U11761 ( .B(n15843), .A(n12631), .S(n13277), .Y(n4592) );
  NAND2X1 U11762 ( .A(n13279), .B(InData[1]), .Y(n12631) );
  INVX1 U11763 ( .A(N3814), .Y(n15843) );
  OAI21X1 U11764 ( .A(n15844), .B(n13277), .C(n13278), .Y(n4591) );
  NAND2X1 U11765 ( .A(n13277), .B(n12630), .Y(n13278) );
  INVX1 U11766 ( .A(N3818), .Y(n15844) );
  MUX2X1 U11767 ( .B(n15845), .A(n12621), .S(n13277), .Y(n4590) );
  AND2X1 U11768 ( .A(n12699), .B(n12636), .Y(n13277) );
  INVX1 U11769 ( .A(n13220), .Y(n12636) );
  OAI21X1 U11770 ( .A(n12630), .B(n13280), .C(rst_b), .Y(n13220) );
  NOR2X1 U11771 ( .A(n13281), .B(n13282), .Y(n13280) );
  AND2X1 U11772 ( .A(n13283), .B(n13284), .Y(n12630) );
  OAI21X1 U11773 ( .A(n13191), .B(n13192), .C(n13285), .Y(n13284) );
  NAND2X1 U11774 ( .A(n13279), .B(InData[0]), .Y(n12621) );
  INVX1 U11775 ( .A(n13282), .Y(n13279) );
  NAND3X1 U11776 ( .A(n13285), .B(n13191), .C(dWriteReg[1]), .Y(n13282) );
  INVX1 U11777 ( .A(N3817), .Y(n15845) );
  MUX2X1 U11778 ( .B(n13286), .A(n13287), .S(n13288), .Y(n4589) );
  NOR2X1 U11779 ( .A(n13289), .B(n12680), .Y(n13288) );
  OAI22X1 U11780 ( .A(n13165), .B(n13290), .C(n13291), .D(n13292), .Y(n13287)
         );
  NAND2X1 U11781 ( .A(n13215), .B(N2880), .Y(n13292) );
  OAI21X1 U11782 ( .A(n13293), .B(n13294), .C(n13295), .Y(n13291) );
  NAND2X1 U11783 ( .A(n13296), .B(n13297), .Y(n13295) );
  MUX2X1 U11784 ( .B(n13298), .A(n13299), .S(n12901), .Y(n13297) );
  AOI21X1 U11785 ( .A(\regZ[8][0] ), .B(n12609), .C(n13300), .Y(n13299) );
  NAND3X1 U11786 ( .A(n13301), .B(n13302), .C(n13303), .Y(n13298) );
  NOR2X1 U11787 ( .A(n13304), .B(n13305), .Y(n13303) );
  OAI21X1 U11788 ( .A(n13306), .B(n13307), .C(n13308), .Y(n13305) );
  MUX2X1 U11789 ( .B(n13309), .A(n13310), .S(n12820), .Y(n13308) );
  AND2X1 U11790 ( .A(n13311), .B(n12609), .Y(n13309) );
  INVX1 U11791 ( .A(n13312), .Y(n13306) );
  INVX1 U11792 ( .A(n13313), .Y(n13304) );
  AOI22X1 U11793 ( .A(n13314), .B(n12700), .C(n13315), .D(n12711), .Y(n13313)
         );
  AOI21X1 U11794 ( .A(n12722), .B(n13316), .C(n13317), .Y(n13302) );
  OAI21X1 U11795 ( .A(n13318), .B(n12620), .C(n13319), .Y(n13317) );
  NAND3X1 U11796 ( .A(n13320), .B(n13321), .C(n13322), .Y(n13319) );
  NOR2X1 U11797 ( .A(n13323), .B(n13324), .Y(n13322) );
  INVX1 U11798 ( .A(n13325), .Y(n13324) );
  AOI22X1 U11799 ( .A(n12722), .B(\regZ[19][0] ), .C(n12757), .D(\regZ[23][0] ), .Y(n13325) );
  OAI21X1 U11800 ( .A(n13326), .B(n13327), .C(n13328), .Y(n13323) );
  AOI22X1 U11801 ( .A(\regZ[22][0] ), .B(n12831), .C(\regZ[20][0] ), .D(n12734), .Y(n13328) );
  INVX1 U11802 ( .A(\regZ[18][0] ), .Y(n13327) );
  AOI22X1 U11803 ( .A(\regZ[21][0] ), .B(n12746), .C(\regZ[17][0] ), .D(n12700), .Y(n13321) );
  NOR2X1 U11804 ( .A(n13300), .B(n13329), .Y(n13320) );
  MUX2X1 U11805 ( .B(n13330), .A(n13331), .S(n12820), .Y(n13329) );
  INVX1 U11806 ( .A(\regZ[24][0] ), .Y(n13331) );
  NAND2X1 U11807 ( .A(\regZ[16][0] ), .B(n12609), .Y(n13330) );
  INVX1 U11808 ( .A(n13332), .Y(n13318) );
  AOI22X1 U11809 ( .A(n12757), .B(n13333), .C(n12831), .D(n13334), .Y(n13301)
         );
  AOI22X1 U11810 ( .A(n12688), .B(n13335), .C(n12820), .D(n13336), .Y(n13296)
         );
  NAND3X1 U11811 ( .A(n13337), .B(n13338), .C(n13339), .Y(n13336) );
  NOR2X1 U11812 ( .A(n13340), .B(n13341), .Y(n13339) );
  OAI22X1 U11813 ( .A(n13342), .B(n12685), .C(n13343), .D(n13326), .Y(n13341)
         );
  OAI21X1 U11814 ( .A(n13344), .B(n13307), .C(n13345), .Y(n13340) );
  NAND3X1 U11815 ( .A(n12901), .B(n13346), .C(n12609), .Y(n13345) );
  INVX1 U11816 ( .A(n12819), .Y(n12901) );
  AOI22X1 U11817 ( .A(n12757), .B(n13347), .C(n12746), .D(n13348), .Y(n13338)
         );
  AOI22X1 U11818 ( .A(n12700), .B(n13349), .C(n12722), .D(n13350), .Y(n13337)
         );
  NAND3X1 U11819 ( .A(n13351), .B(n13352), .C(n13353), .Y(n13335) );
  NOR2X1 U11820 ( .A(n13354), .B(n13355), .Y(n13353) );
  INVX1 U11821 ( .A(n13356), .Y(n13355) );
  AOI22X1 U11822 ( .A(n13357), .B(n12757), .C(n13358), .D(n12700), .Y(n13356)
         );
  OAI21X1 U11823 ( .A(n13359), .B(n13326), .C(n13300), .Y(n13354) );
  OAI21X1 U11824 ( .A(n13360), .B(n12758), .C(n13361), .Y(n13300) );
  OAI21X1 U11825 ( .A(n13362), .B(n13363), .C(n12820), .Y(n13361) );
  OAI21X1 U11826 ( .A(n13364), .B(n13365), .C(n13366), .Y(n13363) );
  AOI22X1 U11827 ( .A(\regZ[11][0] ), .B(n12722), .C(\regZ[13][0] ), .D(n12746), .Y(n13366) );
  NAND2X1 U11828 ( .A(n13367), .B(n13368), .Y(n13362) );
  AOI22X1 U11829 ( .A(\regZ[14][0] ), .B(n12831), .C(\regZ[12][0] ), .D(n12734), .Y(n13368) );
  INVX1 U11830 ( .A(n12685), .Y(n12831) );
  NAND3X1 U11831 ( .A(n13369), .B(n13370), .C(n13371), .Y(n12685) );
  AOI22X1 U11832 ( .A(\regZ[10][0] ), .B(n12711), .C(\regZ[15][0] ), .D(n12757), .Y(n13367) );
  INVX1 U11833 ( .A(n12688), .Y(n12758) );
  NOR2X1 U11834 ( .A(n13372), .B(n13373), .Y(n13360) );
  OAI21X1 U11835 ( .A(n13374), .B(n13375), .C(n13376), .Y(n13373) );
  AOI22X1 U11836 ( .A(\regZ[5][0] ), .B(n12746), .C(\regZ[1][0] ), .D(n12700), 
        .Y(n13376) );
  INVX1 U11837 ( .A(n13364), .Y(n12700) );
  NAND3X1 U11838 ( .A(n13377), .B(n13378), .C(n13379), .Y(n13364) );
  INVX1 U11839 ( .A(\regZ[0][0] ), .Y(n13375) );
  NAND2X1 U11840 ( .A(n13380), .B(n13381), .Y(n13372) );
  AOI22X1 U11841 ( .A(\regZ[4][0] ), .B(n12734), .C(\regZ[2][0] ), .D(n12711), 
        .Y(n13381) );
  INVX1 U11842 ( .A(n13326), .Y(n12711) );
  AOI22X1 U11843 ( .A(\regZ[7][0] ), .B(n12757), .C(\regZ[3][0] ), .D(n12722), 
        .Y(n13380) );
  INVX1 U11844 ( .A(n12596), .Y(n12757) );
  NAND3X1 U11845 ( .A(n13370), .B(n13378), .C(n13369), .Y(n12596) );
  NAND3X1 U11846 ( .A(n13377), .B(n13370), .C(n13371), .Y(n13326) );
  INVX1 U11847 ( .A(n13382), .Y(n13359) );
  AOI22X1 U11848 ( .A(n12734), .B(n13383), .C(n12722), .D(n13384), .Y(n13352)
         );
  INVX1 U11849 ( .A(n13385), .Y(n12722) );
  NAND3X1 U11850 ( .A(n13370), .B(n13378), .C(n13377), .Y(n13385) );
  INVX1 U11851 ( .A(n13307), .Y(n12734) );
  NAND3X1 U11852 ( .A(n13369), .B(n13379), .C(n13371), .Y(n13307) );
  AOI22X1 U11853 ( .A(n12609), .B(n13386), .C(n12746), .D(n13387), .Y(n13351)
         );
  INVX1 U11854 ( .A(n12620), .Y(n12746) );
  NAND3X1 U11855 ( .A(n13369), .B(n13378), .C(n13379), .Y(n12620) );
  INVX1 U11856 ( .A(n13371), .Y(n13378) );
  INVX1 U11857 ( .A(n13377), .Y(n13369) );
  INVX1 U11858 ( .A(n13374), .Y(n12609) );
  NAND3X1 U11859 ( .A(n13379), .B(n13377), .C(n13371), .Y(n13374) );
  AOI21X1 U11860 ( .A(n13388), .B(n13389), .C(n13390), .Y(n13371) );
  XOR2X1 U11861 ( .A(n13391), .B(n13392), .Y(n13377) );
  XOR2X1 U11862 ( .A(n13393), .B(n13394), .Y(n13391) );
  INVX1 U11863 ( .A(n13370), .Y(n13379) );
  XOR2X1 U11864 ( .A(n13395), .B(n13396), .Y(n13370) );
  XNOR2X1 U11865 ( .A(n13390), .B(n13397), .Y(n13395) );
  NOR2X1 U11866 ( .A(n12820), .B(n12819), .Y(n12688) );
  XNOR2X1 U11867 ( .A(n13398), .B(n13399), .Y(n12819) );
  XOR2X1 U11868 ( .A(n13188), .B(n13187), .Y(n13398) );
  AOI21X1 U11869 ( .A(n13400), .B(n13401), .C(n13402), .Y(n13187) );
  INVX1 U11870 ( .A(n13403), .Y(n13402) );
  OAI21X1 U11871 ( .A(n13401), .B(n13400), .C(n13404), .Y(n13403) );
  OAI21X1 U11872 ( .A(n13405), .B(n13406), .C(n13407), .Y(n13188) );
  INVX1 U11873 ( .A(N3193), .Y(n13406) );
  XOR2X1 U11874 ( .A(n13408), .B(n13401), .Y(n12820) );
  OAI21X1 U11875 ( .A(n13393), .B(n13392), .C(n13409), .Y(n13401) );
  INVX1 U11876 ( .A(n13410), .Y(n13409) );
  AOI21X1 U11877 ( .A(n13393), .B(n13392), .C(n13394), .Y(n13410) );
  AOI22X1 U11878 ( .A(n13411), .B(n15325), .C(n13412), .D(n15327), .Y(n13394)
         );
  OAI21X1 U11879 ( .A(n13405), .B(n13413), .C(n13407), .Y(n13392) );
  INVX1 U11880 ( .A(n13414), .Y(n13407) );
  INVX1 U11881 ( .A(N3191), .Y(n13413) );
  OAI21X1 U11882 ( .A(n13415), .B(n13416), .C(n13417), .Y(n13393) );
  OAI21X1 U11883 ( .A(n13397), .B(n13396), .C(n13390), .Y(n13417) );
  NOR2X1 U11884 ( .A(n13388), .B(n13389), .Y(n13390) );
  AOI22X1 U11885 ( .A(dx[0]), .B(n15325), .C(n15327), .D(N3189), .Y(n13389) );
  INVX1 U11886 ( .A(n13415), .Y(n13396) );
  INVX1 U11887 ( .A(n13416), .Y(n13397) );
  OAI22X1 U11888 ( .A(n13418), .B(n13419), .C(n13420), .D(n13405), .Y(n13416)
         );
  AOI21X1 U11889 ( .A(n15327), .B(N3190), .C(n13414), .Y(n13415) );
  XOR2X1 U11890 ( .A(n13404), .B(n13400), .Y(n13408) );
  OAI21X1 U11891 ( .A(n13421), .B(n13405), .C(n13422), .Y(n13400) );
  AOI21X1 U11892 ( .A(n15327), .B(N3192), .C(n13414), .Y(n13404) );
  NOR2X1 U11893 ( .A(n13419), .B(n12539), .Y(n13414) );
  OAI21X1 U11894 ( .A(n13423), .B(n13424), .C(n13425), .Y(n13294) );
  OAI21X1 U11895 ( .A(n13426), .B(n13427), .C(n13428), .Y(n13425) );
  MUX2X1 U11896 ( .B(n13429), .A(n13430), .S(n13431), .Y(n13427) );
  NOR2X1 U11897 ( .A(n13432), .B(n13433), .Y(n13430) );
  OAI22X1 U11898 ( .A(n13343), .B(n13434), .C(n13344), .D(n13435), .Y(n13433)
         );
  INVX1 U11899 ( .A(n13436), .Y(n13344) );
  NAND3X1 U11900 ( .A(n13437), .B(n13438), .C(n13439), .Y(n13436) );
  NOR2X1 U11901 ( .A(\regZ[12][1] ), .B(n13440), .Y(n13439) );
  OR2X1 U11902 ( .A(\regZ[12][3] ), .B(\regZ[12][2] ), .Y(n13440) );
  NOR2X1 U11903 ( .A(\regZ[12][7] ), .B(\regZ[12][6] ), .Y(n13438) );
  NOR2X1 U11904 ( .A(\regZ[12][5] ), .B(\regZ[12][4] ), .Y(n13437) );
  INVX1 U11905 ( .A(n13441), .Y(n13343) );
  NAND3X1 U11906 ( .A(n13442), .B(n13443), .C(n13444), .Y(n13441) );
  NOR2X1 U11907 ( .A(\regZ[10][1] ), .B(n13445), .Y(n13444) );
  OR2X1 U11908 ( .A(\regZ[10][3] ), .B(\regZ[10][2] ), .Y(n13445) );
  NOR2X1 U11909 ( .A(\regZ[10][7] ), .B(\regZ[10][6] ), .Y(n13443) );
  NOR2X1 U11910 ( .A(\regZ[10][5] ), .B(\regZ[10][4] ), .Y(n13442) );
  OAI21X1 U11911 ( .A(n13342), .B(n13446), .C(n13447), .Y(n13432) );
  NAND3X1 U11912 ( .A(n13448), .B(n13346), .C(n13449), .Y(n13447) );
  NAND3X1 U11913 ( .A(n13450), .B(n13451), .C(n13452), .Y(n13346) );
  NOR2X1 U11914 ( .A(\regZ[8][1] ), .B(n13453), .Y(n13452) );
  OR2X1 U11915 ( .A(\regZ[8][3] ), .B(\regZ[8][2] ), .Y(n13453) );
  NOR2X1 U11916 ( .A(\regZ[8][7] ), .B(\regZ[8][6] ), .Y(n13451) );
  NOR2X1 U11917 ( .A(\regZ[8][5] ), .B(\regZ[8][4] ), .Y(n13450) );
  INVX1 U11918 ( .A(n13454), .Y(n13342) );
  NAND3X1 U11919 ( .A(n13455), .B(n13456), .C(n13457), .Y(n13454) );
  NOR2X1 U11920 ( .A(\regZ[14][1] ), .B(n13458), .Y(n13457) );
  OR2X1 U11921 ( .A(\regZ[14][3] ), .B(\regZ[14][2] ), .Y(n13458) );
  NOR2X1 U11922 ( .A(\regZ[14][7] ), .B(\regZ[14][6] ), .Y(n13456) );
  NOR2X1 U11923 ( .A(\regZ[14][5] ), .B(\regZ[14][4] ), .Y(n13455) );
  AND2X1 U11924 ( .A(n13459), .B(n13460), .Y(n13429) );
  AOI22X1 U11925 ( .A(n13349), .B(n13448), .C(n13350), .D(n13461), .Y(n13460)
         );
  NAND3X1 U11926 ( .A(n13462), .B(n13463), .C(n13464), .Y(n13350) );
  NOR2X1 U11927 ( .A(\regZ[11][1] ), .B(n13465), .Y(n13464) );
  OR2X1 U11928 ( .A(\regZ[11][3] ), .B(\regZ[11][2] ), .Y(n13465) );
  NOR2X1 U11929 ( .A(\regZ[11][7] ), .B(\regZ[11][6] ), .Y(n13463) );
  NOR2X1 U11930 ( .A(\regZ[11][5] ), .B(\regZ[11][4] ), .Y(n13462) );
  NAND3X1 U11931 ( .A(n13466), .B(n13467), .C(n13468), .Y(n13349) );
  NOR2X1 U11932 ( .A(\regZ[9][1] ), .B(n13469), .Y(n13468) );
  OR2X1 U11933 ( .A(\regZ[9][3] ), .B(\regZ[9][2] ), .Y(n13469) );
  NOR2X1 U11934 ( .A(\regZ[9][7] ), .B(\regZ[9][6] ), .Y(n13467) );
  NOR2X1 U11935 ( .A(\regZ[9][5] ), .B(\regZ[9][4] ), .Y(n13466) );
  AOI22X1 U11936 ( .A(n13348), .B(n13470), .C(n13347), .D(n13471), .Y(n13459)
         );
  NAND3X1 U11937 ( .A(n13472), .B(n13473), .C(n13474), .Y(n13347) );
  NOR2X1 U11938 ( .A(\regZ[15][1] ), .B(n13475), .Y(n13474) );
  OR2X1 U11939 ( .A(\regZ[15][3] ), .B(\regZ[15][2] ), .Y(n13475) );
  NOR2X1 U11940 ( .A(\regZ[15][7] ), .B(\regZ[15][6] ), .Y(n13473) );
  NOR2X1 U11941 ( .A(\regZ[15][5] ), .B(\regZ[15][4] ), .Y(n13472) );
  NAND3X1 U11942 ( .A(n13476), .B(n13477), .C(n13478), .Y(n13348) );
  NOR2X1 U11943 ( .A(\regZ[13][1] ), .B(n13479), .Y(n13478) );
  OR2X1 U11944 ( .A(\regZ[13][3] ), .B(\regZ[13][2] ), .Y(n13479) );
  NOR2X1 U11945 ( .A(\regZ[13][7] ), .B(\regZ[13][6] ), .Y(n13477) );
  NOR2X1 U11946 ( .A(\regZ[13][5] ), .B(\regZ[13][4] ), .Y(n13476) );
  AND2X1 U11947 ( .A(n13310), .B(n13480), .Y(n13426) );
  NAND3X1 U11948 ( .A(n13481), .B(n13482), .C(n13483), .Y(n13310) );
  NOR2X1 U11949 ( .A(\regZ[24][1] ), .B(n13484), .Y(n13483) );
  OR2X1 U11950 ( .A(\regZ[24][3] ), .B(\regZ[24][2] ), .Y(n13484) );
  NOR2X1 U11951 ( .A(\regZ[24][7] ), .B(\regZ[24][6] ), .Y(n13482) );
  NOR2X1 U11952 ( .A(\regZ[24][5] ), .B(\regZ[24][4] ), .Y(n13481) );
  NAND2X1 U11953 ( .A(n13485), .B(n13486), .Y(n13424) );
  OAI21X1 U11954 ( .A(n13487), .B(n13488), .C(n13489), .Y(n13486) );
  INVX1 U11955 ( .A(n13490), .Y(n13488) );
  AOI22X1 U11956 ( .A(n13448), .B(\regZ[0][0] ), .C(n13461), .D(\regZ[2][0] ), 
        .Y(n13490) );
  OAI21X1 U11957 ( .A(n13435), .B(n13491), .C(n13492), .Y(n13487) );
  NAND2X1 U11958 ( .A(\regZ[6][0] ), .B(n13471), .Y(n13492) );
  INVX1 U11959 ( .A(\regZ[4][0] ), .Y(n13491) );
  INVX1 U11960 ( .A(n13493), .Y(n13485) );
  AOI21X1 U11961 ( .A(n13494), .B(n13495), .C(n13496), .Y(n13493) );
  AOI22X1 U11962 ( .A(n13448), .B(\regZ[1][0] ), .C(n13461), .D(\regZ[3][0] ), 
        .Y(n13495) );
  AOI22X1 U11963 ( .A(n13470), .B(\regZ[5][0] ), .C(n13471), .D(\regZ[7][0] ), 
        .Y(n13494) );
  OAI21X1 U11964 ( .A(n13497), .B(n13498), .C(n13499), .Y(n13423) );
  OAI21X1 U11965 ( .A(n13500), .B(n13501), .C(n13502), .Y(n13499) );
  OAI21X1 U11966 ( .A(n13449), .B(n13503), .C(n13504), .Y(n13502) );
  OAI21X1 U11967 ( .A(n13446), .B(n13505), .C(n13506), .Y(n13501) );
  OAI21X1 U11968 ( .A(\regZ[24][0] ), .B(n13507), .C(n13480), .Y(n13506) );
  INVX1 U11969 ( .A(n13503), .Y(n13507) );
  MUX2X1 U11970 ( .B(n13508), .A(n13509), .S(n13431), .Y(n13503) );
  NAND2X1 U11971 ( .A(n13510), .B(n13511), .Y(n13509) );
  AOI22X1 U11972 ( .A(n13512), .B(\regZ[16][0] ), .C(\regZ[22][0] ), .D(n13471), .Y(n13511) );
  NOR2X1 U11973 ( .A(n13428), .B(n13513), .Y(n13512) );
  AOI22X1 U11974 ( .A(\regZ[20][0] ), .B(n13470), .C(\regZ[18][0] ), .D(n13461), .Y(n13510) );
  NAND2X1 U11975 ( .A(n13514), .B(n13515), .Y(n13508) );
  AOI22X1 U11976 ( .A(\regZ[23][0] ), .B(n13471), .C(\regZ[21][0] ), .D(n13470), .Y(n13515) );
  AOI22X1 U11977 ( .A(\regZ[19][0] ), .B(n13461), .C(\regZ[17][0] ), .D(n13448), .Y(n13514) );
  MUX2X1 U11978 ( .B(\regZ[15][0] ), .A(\regZ[14][0] ), .S(n13431), .Y(n13505)
         );
  MUX2X1 U11979 ( .B(n13516), .A(n13517), .S(n13431), .Y(n13500) );
  AOI22X1 U11980 ( .A(\regZ[12][0] ), .B(n13470), .C(\regZ[10][0] ), .D(n13461), .Y(n13517) );
  INVX1 U11981 ( .A(n13518), .Y(n13516) );
  OAI21X1 U11982 ( .A(n13365), .B(n13513), .C(n13519), .Y(n13518) );
  AOI22X1 U11983 ( .A(n13461), .B(\regZ[11][0] ), .C(n13470), .D(\regZ[13][0] ), .Y(n13519) );
  INVX1 U11984 ( .A(\regZ[9][0] ), .Y(n13365) );
  NAND2X1 U11985 ( .A(n13428), .B(\regZ[8][0] ), .Y(n13498) );
  INVX1 U11986 ( .A(n13504), .Y(n13428) );
  NAND3X1 U11987 ( .A(n13448), .B(n13431), .C(n13449), .Y(n13497) );
  NAND3X1 U11988 ( .A(n13520), .B(n13521), .C(n13522), .Y(n13293) );
  INVX1 U11989 ( .A(n13523), .Y(n13522) );
  AOI21X1 U11990 ( .A(n13524), .B(n13525), .C(n13496), .Y(n13523) );
  NAND3X1 U11991 ( .A(n13526), .B(n13504), .C(n13449), .Y(n13496) );
  INVX1 U11992 ( .A(n13431), .Y(n13526) );
  AOI22X1 U11993 ( .A(n13358), .B(n13448), .C(n13384), .D(n13461), .Y(n13525)
         );
  NAND3X1 U11994 ( .A(n13527), .B(n13528), .C(n13529), .Y(n13384) );
  NOR2X1 U11995 ( .A(\regZ[3][1] ), .B(n13530), .Y(n13529) );
  OR2X1 U11996 ( .A(\regZ[3][3] ), .B(\regZ[3][2] ), .Y(n13530) );
  NOR2X1 U11997 ( .A(\regZ[3][7] ), .B(\regZ[3][6] ), .Y(n13528) );
  NOR2X1 U11998 ( .A(\regZ[3][5] ), .B(\regZ[3][4] ), .Y(n13527) );
  NAND3X1 U11999 ( .A(n13531), .B(n13532), .C(n13533), .Y(n13358) );
  NOR2X1 U12000 ( .A(\regZ[1][1] ), .B(n13534), .Y(n13533) );
  OR2X1 U12001 ( .A(\regZ[1][3] ), .B(\regZ[1][2] ), .Y(n13534) );
  NOR2X1 U12002 ( .A(\regZ[1][7] ), .B(\regZ[1][6] ), .Y(n13532) );
  NOR2X1 U12003 ( .A(\regZ[1][5] ), .B(\regZ[1][4] ), .Y(n13531) );
  AOI22X1 U12004 ( .A(n13387), .B(n13470), .C(n13357), .D(n13471), .Y(n13524)
         );
  NAND3X1 U12005 ( .A(n13535), .B(n13536), .C(n13537), .Y(n13357) );
  NOR2X1 U12006 ( .A(\regZ[7][1] ), .B(n13538), .Y(n13537) );
  OR2X1 U12007 ( .A(\regZ[7][3] ), .B(\regZ[7][2] ), .Y(n13538) );
  NOR2X1 U12008 ( .A(\regZ[7][7] ), .B(\regZ[7][6] ), .Y(n13536) );
  NOR2X1 U12009 ( .A(\regZ[7][5] ), .B(\regZ[7][4] ), .Y(n13535) );
  NAND3X1 U12010 ( .A(n13539), .B(n13540), .C(n13541), .Y(n13387) );
  NOR2X1 U12011 ( .A(\regZ[5][1] ), .B(n13542), .Y(n13541) );
  OR2X1 U12012 ( .A(\regZ[5][3] ), .B(\regZ[5][2] ), .Y(n13542) );
  NOR2X1 U12013 ( .A(\regZ[5][7] ), .B(\regZ[5][6] ), .Y(n13540) );
  NOR2X1 U12014 ( .A(\regZ[5][5] ), .B(\regZ[5][4] ), .Y(n13539) );
  NAND2X1 U12015 ( .A(n13543), .B(n13480), .Y(n13521) );
  MUX2X1 U12016 ( .B(n13544), .A(n13545), .S(n13431), .Y(n13543) );
  NOR2X1 U12017 ( .A(n13546), .B(n13547), .Y(n13545) );
  INVX1 U12018 ( .A(n13548), .Y(n13547) );
  AOI22X1 U12019 ( .A(n13315), .B(n13461), .C(n13312), .D(n13470), .Y(n13548)
         );
  NAND3X1 U12020 ( .A(n13549), .B(n13550), .C(n13551), .Y(n13312) );
  NOR2X1 U12021 ( .A(\regZ[20][1] ), .B(n13552), .Y(n13551) );
  OR2X1 U12022 ( .A(\regZ[20][3] ), .B(\regZ[20][2] ), .Y(n13552) );
  NOR2X1 U12023 ( .A(\regZ[20][7] ), .B(\regZ[20][6] ), .Y(n13550) );
  NOR2X1 U12024 ( .A(\regZ[20][5] ), .B(\regZ[20][4] ), .Y(n13549) );
  NAND3X1 U12025 ( .A(n13553), .B(n13554), .C(n13555), .Y(n13315) );
  NOR2X1 U12026 ( .A(\regZ[18][1] ), .B(n13556), .Y(n13555) );
  OR2X1 U12027 ( .A(\regZ[18][3] ), .B(\regZ[18][2] ), .Y(n13556) );
  NOR2X1 U12028 ( .A(\regZ[18][7] ), .B(\regZ[18][6] ), .Y(n13554) );
  NOR2X1 U12029 ( .A(\regZ[18][5] ), .B(\regZ[18][4] ), .Y(n13553) );
  OAI21X1 U12030 ( .A(n13557), .B(n13446), .C(n13558), .Y(n13546) );
  NAND3X1 U12031 ( .A(n13504), .B(n13311), .C(n13448), .Y(n13558) );
  NAND3X1 U12032 ( .A(n13559), .B(n13560), .C(n13561), .Y(n13311) );
  NOR2X1 U12033 ( .A(\regZ[16][1] ), .B(n13562), .Y(n13561) );
  OR2X1 U12034 ( .A(\regZ[16][3] ), .B(\regZ[16][2] ), .Y(n13562) );
  NOR2X1 U12035 ( .A(\regZ[16][7] ), .B(\regZ[16][6] ), .Y(n13560) );
  NOR2X1 U12036 ( .A(\regZ[16][5] ), .B(\regZ[16][4] ), .Y(n13559) );
  INVX1 U12037 ( .A(n13471), .Y(n13446) );
  INVX1 U12038 ( .A(n13334), .Y(n13557) );
  NAND3X1 U12039 ( .A(n13563), .B(n13564), .C(n13565), .Y(n13334) );
  NOR2X1 U12040 ( .A(\regZ[22][1] ), .B(n13566), .Y(n13565) );
  OR2X1 U12041 ( .A(\regZ[22][3] ), .B(\regZ[22][2] ), .Y(n13566) );
  NOR2X1 U12042 ( .A(\regZ[22][7] ), .B(\regZ[22][6] ), .Y(n13564) );
  NOR2X1 U12043 ( .A(\regZ[22][5] ), .B(\regZ[22][4] ), .Y(n13563) );
  AND2X1 U12044 ( .A(n13567), .B(n13568), .Y(n13544) );
  AOI22X1 U12045 ( .A(n13314), .B(n13448), .C(n13316), .D(n13461), .Y(n13568)
         );
  NAND3X1 U12046 ( .A(n13569), .B(n13570), .C(n13571), .Y(n13316) );
  NOR2X1 U12047 ( .A(\regZ[19][1] ), .B(n13572), .Y(n13571) );
  OR2X1 U12048 ( .A(\regZ[19][3] ), .B(\regZ[19][2] ), .Y(n13572) );
  NOR2X1 U12049 ( .A(\regZ[19][7] ), .B(\regZ[19][6] ), .Y(n13570) );
  NOR2X1 U12050 ( .A(\regZ[19][5] ), .B(\regZ[19][4] ), .Y(n13569) );
  NAND3X1 U12051 ( .A(n13573), .B(n13574), .C(n13575), .Y(n13314) );
  NOR2X1 U12052 ( .A(\regZ[17][1] ), .B(n13576), .Y(n13575) );
  OR2X1 U12053 ( .A(\regZ[17][3] ), .B(\regZ[17][2] ), .Y(n13576) );
  NOR2X1 U12054 ( .A(\regZ[17][7] ), .B(\regZ[17][6] ), .Y(n13574) );
  NOR2X1 U12055 ( .A(\regZ[17][5] ), .B(\regZ[17][4] ), .Y(n13573) );
  AOI22X1 U12056 ( .A(n13332), .B(n13470), .C(n13333), .D(n13471), .Y(n13567)
         );
  NAND3X1 U12057 ( .A(n13577), .B(n13578), .C(n13579), .Y(n13333) );
  NOR2X1 U12058 ( .A(\regZ[23][1] ), .B(n13580), .Y(n13579) );
  OR2X1 U12059 ( .A(\regZ[23][3] ), .B(\regZ[23][2] ), .Y(n13580) );
  NOR2X1 U12060 ( .A(\regZ[23][7] ), .B(\regZ[23][6] ), .Y(n13578) );
  NOR2X1 U12061 ( .A(\regZ[23][5] ), .B(\regZ[23][4] ), .Y(n13577) );
  NAND3X1 U12062 ( .A(n13581), .B(n13582), .C(n13583), .Y(n13332) );
  NOR2X1 U12063 ( .A(\regZ[21][1] ), .B(n13584), .Y(n13583) );
  OR2X1 U12064 ( .A(\regZ[21][3] ), .B(\regZ[21][2] ), .Y(n13584) );
  NOR2X1 U12065 ( .A(\regZ[21][7] ), .B(\regZ[21][6] ), .Y(n13582) );
  NOR2X1 U12066 ( .A(\regZ[21][5] ), .B(\regZ[21][4] ), .Y(n13581) );
  OAI21X1 U12067 ( .A(n13585), .B(n13586), .C(n13489), .Y(n13520) );
  INVX1 U12068 ( .A(n13587), .Y(n13489) );
  NAND3X1 U12069 ( .A(n13504), .B(n13431), .C(n13449), .Y(n13587) );
  INVX1 U12070 ( .A(n13480), .Y(n13449) );
  XNOR2X1 U12071 ( .A(n13588), .B(n13589), .Y(n13480) );
  XNOR2X1 U12072 ( .A(dx[1]), .B(n13590), .Y(n13589) );
  XOR2X1 U12073 ( .A(n13591), .B(n13592), .Y(n13588) );
  NOR2X1 U12074 ( .A(n13593), .B(n13594), .Y(n13592) );
  INVX1 U12075 ( .A(n13595), .Y(n13593) );
  OAI21X1 U12076 ( .A(n13596), .B(n13421), .C(n13597), .Y(n13591) );
  OAI21X1 U12077 ( .A(n13598), .B(n13599), .C(dx[1]), .Y(n13597) );
  INVX1 U12078 ( .A(n13421), .Y(n13598) );
  OAI21X1 U12079 ( .A(dx[0]), .B(n13388), .C(n13600), .Y(n13431) );
  XOR2X1 U12080 ( .A(n13601), .B(n13421), .Y(n13504) );
  XOR2X1 U12081 ( .A(n13594), .B(n13595), .Y(n13421) );
  XOR2X1 U12082 ( .A(n13602), .B(n13405), .Y(n13594) );
  XNOR2X1 U12083 ( .A(n13596), .B(dx[1]), .Y(n13601) );
  INVX1 U12084 ( .A(n13599), .Y(n13596) );
  OAI21X1 U12085 ( .A(n13603), .B(n13604), .C(n13605), .Y(n13599) );
  OAI21X1 U12086 ( .A(n13606), .B(n13412), .C(dx[1]), .Y(n13605) );
  INVX1 U12087 ( .A(n13604), .Y(n13606) );
  INVX1 U12088 ( .A(n13607), .Y(n13586) );
  AOI22X1 U12089 ( .A(n13386), .B(n13448), .C(n13382), .D(n13461), .Y(n13607)
         );
  INVX1 U12090 ( .A(n13434), .Y(n13461) );
  NAND2X1 U12091 ( .A(n13608), .B(n13609), .Y(n13434) );
  NAND3X1 U12092 ( .A(n13610), .B(n13611), .C(n13612), .Y(n13382) );
  NOR2X1 U12093 ( .A(\regZ[2][1] ), .B(n13613), .Y(n13612) );
  OR2X1 U12094 ( .A(\regZ[2][3] ), .B(\regZ[2][2] ), .Y(n13613) );
  NOR2X1 U12095 ( .A(\regZ[2][7] ), .B(\regZ[2][6] ), .Y(n13611) );
  NOR2X1 U12096 ( .A(\regZ[2][5] ), .B(\regZ[2][4] ), .Y(n13610) );
  INVX1 U12097 ( .A(n13513), .Y(n13448) );
  NAND2X1 U12098 ( .A(n13614), .B(n13609), .Y(n13513) );
  NAND3X1 U12099 ( .A(n13615), .B(n13616), .C(n13617), .Y(n13386) );
  NOR2X1 U12100 ( .A(\regZ[0][1] ), .B(n13618), .Y(n13617) );
  OR2X1 U12101 ( .A(\regZ[0][3] ), .B(\regZ[0][2] ), .Y(n13618) );
  NOR2X1 U12102 ( .A(\regZ[0][7] ), .B(\regZ[0][6] ), .Y(n13616) );
  NOR2X1 U12103 ( .A(\regZ[0][5] ), .B(\regZ[0][4] ), .Y(n13615) );
  OAI21X1 U12104 ( .A(n13619), .B(n13435), .C(n13620), .Y(n13585) );
  OAI21X1 U12105 ( .A(n13621), .B(n13622), .C(n13471), .Y(n13620) );
  NOR2X1 U12106 ( .A(n13609), .B(n13614), .Y(n13471) );
  OR2X1 U12107 ( .A(\regZ[6][1] ), .B(n13623), .Y(n13622) );
  OR2X1 U12108 ( .A(\regZ[6][3] ), .B(\regZ[6][2] ), .Y(n13623) );
  NAND2X1 U12109 ( .A(n13624), .B(n13625), .Y(n13621) );
  NOR2X1 U12110 ( .A(\regZ[6][7] ), .B(\regZ[6][6] ), .Y(n13625) );
  NOR2X1 U12111 ( .A(\regZ[6][5] ), .B(\regZ[6][4] ), .Y(n13624) );
  INVX1 U12112 ( .A(n13470), .Y(n13435) );
  NOR2X1 U12113 ( .A(n13609), .B(n13608), .Y(n13470) );
  INVX1 U12114 ( .A(n13614), .Y(n13608) );
  XOR2X1 U12115 ( .A(n13420), .B(n13626), .Y(n13614) );
  XNOR2X1 U12116 ( .A(n12539), .B(n13627), .Y(n13626) );
  XOR2X1 U12117 ( .A(n13628), .B(n13604), .Y(n13609) );
  OAI21X1 U12118 ( .A(n13627), .B(n13629), .C(n13630), .Y(n13604) );
  OAI21X1 U12119 ( .A(n13420), .B(n13600), .C(n12539), .Y(n13630) );
  INVX1 U12120 ( .A(dx[1]), .Y(n12539) );
  INVX1 U12121 ( .A(n13627), .Y(n13600) );
  INVX1 U12122 ( .A(n13420), .Y(n13629) );
  AOI21X1 U12123 ( .A(n13631), .B(n13632), .C(n13633), .Y(n13420) );
  NOR2X1 U12124 ( .A(n13634), .B(n13631), .Y(n13627) );
  XNOR2X1 U12125 ( .A(dx[1]), .B(n13603), .Y(n13628) );
  INVX1 U12126 ( .A(n13412), .Y(n13603) );
  OAI21X1 U12127 ( .A(n13633), .B(n13635), .C(n13595), .Y(n13412) );
  NAND2X1 U12128 ( .A(n13633), .B(n13635), .Y(n13595) );
  XNOR2X1 U12129 ( .A(n13636), .B(n15327), .Y(n13635) );
  MUX2X1 U12130 ( .B(n13637), .A(n13638), .S(n13405), .Y(n13633) );
  INVX1 U12131 ( .A(n13383), .Y(n13619) );
  NAND3X1 U12132 ( .A(n13639), .B(n13640), .C(n13641), .Y(n13383) );
  NOR2X1 U12133 ( .A(\regZ[4][1] ), .B(n13642), .Y(n13641) );
  OR2X1 U12134 ( .A(\regZ[4][3] ), .B(\regZ[4][2] ), .Y(n13642) );
  NOR2X1 U12135 ( .A(\regZ[4][7] ), .B(\regZ[4][6] ), .Y(n13640) );
  NOR2X1 U12136 ( .A(\regZ[4][5] ), .B(\regZ[4][4] ), .Y(n13639) );
  INVX1 U12137 ( .A(N3336), .Y(n13290) );
  INVX1 U12138 ( .A(\Out_bThres[0] ), .Y(n13286) );
  OAI21X1 U12139 ( .A(n13643), .B(n12519), .C(n13644), .Y(n4588) );
  NAND2X1 U12140 ( .A(N2048), .B(n13645), .Y(n13644) );
  INVX1 U12141 ( .A(tpSum[7]), .Y(n12519) );
  OAI21X1 U12142 ( .A(n13643), .B(n12522), .C(n13646), .Y(n4587) );
  NAND2X1 U12143 ( .A(N2049), .B(n13645), .Y(n13646) );
  INVX1 U12144 ( .A(tpSum[8]), .Y(n12522) );
  OAI21X1 U12145 ( .A(n13643), .B(n12524), .C(n13647), .Y(n4586) );
  NAND2X1 U12146 ( .A(N2050), .B(n13645), .Y(n13647) );
  INVX1 U12147 ( .A(tpSum[9]), .Y(n12524) );
  OAI21X1 U12148 ( .A(n13643), .B(n12526), .C(n13648), .Y(n4585) );
  NAND2X1 U12149 ( .A(N2051), .B(n13645), .Y(n13648) );
  INVX1 U12150 ( .A(tpSum[10]), .Y(n12526) );
  OAI21X1 U12151 ( .A(n13643), .B(n12528), .C(n13649), .Y(n4584) );
  NAND2X1 U12152 ( .A(N2052), .B(n13645), .Y(n13649) );
  INVX1 U12153 ( .A(tpSum[11]), .Y(n12528) );
  OAI21X1 U12154 ( .A(n13643), .B(n12530), .C(n13650), .Y(n4583) );
  NAND2X1 U12155 ( .A(N2053), .B(n13645), .Y(n13650) );
  INVX1 U12156 ( .A(tpSum[12]), .Y(n12530) );
  OAI21X1 U12157 ( .A(n13643), .B(n12532), .C(n13651), .Y(n4582) );
  NAND2X1 U12158 ( .A(N2054), .B(n13645), .Y(n13651) );
  INVX1 U12159 ( .A(tpSum[13]), .Y(n12532) );
  OAI21X1 U12160 ( .A(n13643), .B(n12534), .C(n13652), .Y(n4581) );
  NAND2X1 U12161 ( .A(N2055), .B(n13645), .Y(n13652) );
  NOR2X1 U12162 ( .A(n12535), .B(n12462), .Y(n13645) );
  INVX1 U12163 ( .A(tpSum[14]), .Y(n12534) );
  NOR2X1 U12164 ( .A(n12535), .B(n12537), .Y(n13643) );
  NAND3X1 U12165 ( .A(n13653), .B(n12646), .C(n12668), .Y(n12535) );
  OAI21X1 U12166 ( .A(n12533), .B(n13654), .C(n13655), .Y(n4579) );
  MUX2X1 U12167 ( .B(n13656), .A(N4468), .S(n13657), .Y(n13655) );
  OAI21X1 U12168 ( .A(n13658), .B(n13659), .C(n13660), .Y(n13656) );
  AOI22X1 U12169 ( .A(n13661), .B(n13662), .C(Out_gradient[7]), .D(n13663), 
        .Y(n13660) );
  NAND3X1 U12170 ( .A(n13664), .B(n13665), .C(n13666), .Y(n13662) );
  NOR2X1 U12171 ( .A(n13667), .B(n13668), .Y(n13666) );
  OR2X1 U12172 ( .A(n13669), .B(n13670), .Y(n13668) );
  OAI21X1 U12173 ( .A(n13256), .B(n12850), .C(n13671), .Y(n13670) );
  AOI22X1 U12174 ( .A(N1382), .B(n12710), .C(\regX[19][7] ), .D(n13185), .Y(
        n13671) );
  OAI21X1 U12175 ( .A(n12723), .B(n12720), .C(n13672), .Y(n13669) );
  AOI22X1 U12176 ( .A(\regX[5][7] ), .B(n12745), .C(\regX[0][7] ), .D(n12607), 
        .Y(n13672) );
  NAND3X1 U12177 ( .A(n13673), .B(n13674), .C(n13675), .Y(n13667) );
  AOI21X1 U12178 ( .A(\regX[1][7] ), .B(n12699), .C(n13676), .Y(n13675) );
  OAI22X1 U12179 ( .A(n13271), .B(n13174), .C(n13268), .D(n12899), .Y(n13676)
         );
  AOI22X1 U12180 ( .A(\regX[9][7] ), .B(n12781), .C(\regX[8][7] ), .D(n12769), 
        .Y(n13674) );
  AOI22X1 U12181 ( .A(N1622), .B(n12890), .C(N1684), .D(n12632), .Y(n13673) );
  NOR2X1 U12182 ( .A(n13677), .B(n13678), .Y(n13665) );
  OAI21X1 U12183 ( .A(n12735), .B(n12732), .C(n13679), .Y(n13678) );
  AOI22X1 U12184 ( .A(\regX[20][7] ), .B(n12870), .C(\regX[24][7] ), .D(n12817), .Y(n13679) );
  OAI21X1 U12185 ( .A(n13253), .B(n12840), .C(n13680), .Y(n13677) );
  AOI22X1 U12186 ( .A(\regX[7][7] ), .B(n12756), .C(\regX[16][7] ), .D(n12791), 
        .Y(n13680) );
  NOR2X1 U12187 ( .A(n13681), .B(n13682), .Y(n13664) );
  OAI21X1 U12188 ( .A(n12678), .B(n12677), .C(n13683), .Y(n13682) );
  AOI22X1 U12189 ( .A(\regX[15][7] ), .B(n13250), .C(\regX[21][7] ), .D(n12880), .Y(n13683) );
  OAI21X1 U12190 ( .A(n13247), .B(n12829), .C(n13684), .Y(n13681) );
  AOI22X1 U12191 ( .A(\regX[13][7] ), .B(n13259), .C(\regX[17][7] ), .D(n12803), .Y(n13684) );
  INVX1 U12192 ( .A(Out_direction[7]), .Y(n13659) );
  INVX1 U12193 ( .A(Out_gf[7]), .Y(n12533) );
  OAI21X1 U12194 ( .A(n12531), .B(n13654), .C(n13685), .Y(n4577) );
  MUX2X1 U12195 ( .B(n13686), .A(N4471), .S(n13657), .Y(n13685) );
  OAI21X1 U12196 ( .A(n13658), .B(n13687), .C(n13688), .Y(n13686) );
  AOI22X1 U12197 ( .A(n13661), .B(n13689), .C(Out_gradient[6]), .D(n13663), 
        .Y(n13688) );
  NAND3X1 U12198 ( .A(n13690), .B(n13691), .C(n13692), .Y(n13689) );
  NOR2X1 U12199 ( .A(n13693), .B(n13694), .Y(n13692) );
  OR2X1 U12200 ( .A(n13695), .B(n13696), .Y(n13694) );
  OAI21X1 U12201 ( .A(n13256), .B(n12849), .C(n13697), .Y(n13696) );
  AOI22X1 U12202 ( .A(N1381), .B(n12710), .C(\regX[19][6] ), .D(n13185), .Y(
        n13697) );
  OAI21X1 U12203 ( .A(n12723), .B(n12719), .C(n13698), .Y(n13695) );
  AOI22X1 U12204 ( .A(\regX[5][6] ), .B(n12745), .C(\regX[0][6] ), .D(n12607), 
        .Y(n13698) );
  NAND3X1 U12205 ( .A(n13699), .B(n13700), .C(n13701), .Y(n13693) );
  AOI21X1 U12206 ( .A(\regX[1][6] ), .B(n12699), .C(n13702), .Y(n13701) );
  OAI22X1 U12207 ( .A(n13271), .B(n13173), .C(n13268), .D(n12898), .Y(n13702)
         );
  AOI22X1 U12208 ( .A(\regX[9][6] ), .B(n12781), .C(\regX[8][6] ), .D(n12769), 
        .Y(n13700) );
  AOI22X1 U12209 ( .A(N1621), .B(n12890), .C(N1683), .D(n12632), .Y(n13699) );
  NOR2X1 U12210 ( .A(n13703), .B(n13704), .Y(n13691) );
  OAI21X1 U12211 ( .A(n12735), .B(n12731), .C(n13705), .Y(n13704) );
  AOI22X1 U12212 ( .A(\regX[20][6] ), .B(n12870), .C(\regX[24][6] ), .D(n12817), .Y(n13705) );
  OAI21X1 U12213 ( .A(n13253), .B(n12839), .C(n13706), .Y(n13703) );
  AOI22X1 U12214 ( .A(\regX[7][6] ), .B(n12756), .C(\regX[16][6] ), .D(n12791), 
        .Y(n13706) );
  NOR2X1 U12215 ( .A(n13707), .B(n13708), .Y(n13690) );
  OAI21X1 U12216 ( .A(n12678), .B(n12676), .C(n13709), .Y(n13708) );
  AOI22X1 U12217 ( .A(\regX[15][6] ), .B(n13250), .C(\regX[21][6] ), .D(n12880), .Y(n13709) );
  OAI21X1 U12218 ( .A(n13247), .B(n12828), .C(n13710), .Y(n13707) );
  AOI22X1 U12219 ( .A(\regX[13][6] ), .B(n13259), .C(\regX[17][6] ), .D(n12803), .Y(n13710) );
  INVX1 U12220 ( .A(Out_direction[6]), .Y(n13687) );
  INVX1 U12221 ( .A(Out_gf[6]), .Y(n12531) );
  OAI21X1 U12222 ( .A(n12529), .B(n13654), .C(n13711), .Y(n4575) );
  MUX2X1 U12223 ( .B(n13712), .A(N4474), .S(n13657), .Y(n13711) );
  OAI21X1 U12224 ( .A(n13658), .B(n13713), .C(n13714), .Y(n13712) );
  AOI22X1 U12225 ( .A(n13661), .B(n13715), .C(Out_gradient[5]), .D(n13663), 
        .Y(n13714) );
  NAND3X1 U12226 ( .A(n13716), .B(n13717), .C(n13718), .Y(n13715) );
  NOR2X1 U12227 ( .A(n13719), .B(n13720), .Y(n13718) );
  OR2X1 U12228 ( .A(n13721), .B(n13722), .Y(n13720) );
  OAI21X1 U12229 ( .A(n13256), .B(n12848), .C(n13723), .Y(n13722) );
  AOI22X1 U12230 ( .A(N1380), .B(n12710), .C(\regX[19][5] ), .D(n13185), .Y(
        n13723) );
  OAI21X1 U12231 ( .A(n12723), .B(n12718), .C(n13724), .Y(n13721) );
  AOI22X1 U12232 ( .A(\regX[5][5] ), .B(n12745), .C(\regX[0][5] ), .D(n12607), 
        .Y(n13724) );
  NAND3X1 U12233 ( .A(n13725), .B(n13726), .C(n13727), .Y(n13719) );
  AOI21X1 U12234 ( .A(\regX[1][5] ), .B(n12699), .C(n13728), .Y(n13727) );
  OAI22X1 U12235 ( .A(n13271), .B(n13172), .C(n13268), .D(n12897), .Y(n13728)
         );
  AOI22X1 U12236 ( .A(\regX[9][5] ), .B(n12781), .C(\regX[8][5] ), .D(n12769), 
        .Y(n13726) );
  AOI22X1 U12237 ( .A(N1620), .B(n12890), .C(N1682), .D(n12632), .Y(n13725) );
  NOR2X1 U12238 ( .A(n13729), .B(n13730), .Y(n13717) );
  OAI21X1 U12239 ( .A(n12735), .B(n12730), .C(n13731), .Y(n13730) );
  AOI22X1 U12240 ( .A(\regX[20][5] ), .B(n12870), .C(\regX[24][5] ), .D(n12817), .Y(n13731) );
  OAI21X1 U12241 ( .A(n13253), .B(n12838), .C(n13732), .Y(n13729) );
  AOI22X1 U12242 ( .A(\regX[7][5] ), .B(n12756), .C(\regX[16][5] ), .D(n12791), 
        .Y(n13732) );
  NOR2X1 U12243 ( .A(n13733), .B(n13734), .Y(n13716) );
  OAI21X1 U12244 ( .A(n12678), .B(n12675), .C(n13735), .Y(n13734) );
  AOI22X1 U12245 ( .A(\regX[15][5] ), .B(n13250), .C(\regX[21][5] ), .D(n12880), .Y(n13735) );
  OAI21X1 U12246 ( .A(n13247), .B(n12827), .C(n13736), .Y(n13733) );
  AOI22X1 U12247 ( .A(\regX[13][5] ), .B(n13259), .C(\regX[17][5] ), .D(n12803), .Y(n13736) );
  INVX1 U12248 ( .A(Out_direction[5]), .Y(n13713) );
  INVX1 U12249 ( .A(Out_gf[5]), .Y(n12529) );
  OAI21X1 U12250 ( .A(n12527), .B(n13654), .C(n13737), .Y(n4573) );
  MUX2X1 U12251 ( .B(n13738), .A(N4477), .S(n13657), .Y(n13737) );
  OAI21X1 U12252 ( .A(n13658), .B(n13739), .C(n13740), .Y(n13738) );
  AOI22X1 U12253 ( .A(n13661), .B(n13741), .C(Out_gradient[4]), .D(n13663), 
        .Y(n13740) );
  NAND3X1 U12254 ( .A(n13742), .B(n13743), .C(n13744), .Y(n13741) );
  NOR2X1 U12255 ( .A(n13745), .B(n13746), .Y(n13744) );
  OR2X1 U12256 ( .A(n13747), .B(n13748), .Y(n13746) );
  OAI21X1 U12257 ( .A(n13256), .B(n12847), .C(n13749), .Y(n13748) );
  AOI22X1 U12258 ( .A(N1379), .B(n12710), .C(\regX[19][4] ), .D(n13185), .Y(
        n13749) );
  OAI21X1 U12259 ( .A(n12723), .B(n12717), .C(n13750), .Y(n13747) );
  AOI22X1 U12260 ( .A(\regX[5][4] ), .B(n12745), .C(\regX[0][4] ), .D(n12607), 
        .Y(n13750) );
  NAND3X1 U12261 ( .A(n13751), .B(n13752), .C(n13753), .Y(n13745) );
  AOI21X1 U12262 ( .A(\regX[1][4] ), .B(n12699), .C(n13754), .Y(n13753) );
  OAI22X1 U12263 ( .A(n13271), .B(n13171), .C(n13268), .D(n12896), .Y(n13754)
         );
  AOI22X1 U12264 ( .A(\regX[9][4] ), .B(n12781), .C(\regX[8][4] ), .D(n12769), 
        .Y(n13752) );
  AOI22X1 U12265 ( .A(N1619), .B(n12890), .C(N1681), .D(n12632), .Y(n13751) );
  NOR2X1 U12266 ( .A(n13755), .B(n13756), .Y(n13743) );
  OAI21X1 U12267 ( .A(n12735), .B(n12729), .C(n13757), .Y(n13756) );
  AOI22X1 U12268 ( .A(\regX[20][4] ), .B(n12870), .C(\regX[24][4] ), .D(n12817), .Y(n13757) );
  OAI21X1 U12269 ( .A(n13253), .B(n12837), .C(n13758), .Y(n13755) );
  AOI22X1 U12270 ( .A(\regX[7][4] ), .B(n12756), .C(\regX[16][4] ), .D(n12791), 
        .Y(n13758) );
  NOR2X1 U12271 ( .A(n13759), .B(n13760), .Y(n13742) );
  OAI21X1 U12272 ( .A(n12678), .B(n12674), .C(n13761), .Y(n13760) );
  AOI22X1 U12273 ( .A(\regX[15][4] ), .B(n13250), .C(\regX[21][4] ), .D(n12880), .Y(n13761) );
  OAI21X1 U12274 ( .A(n13247), .B(n12826), .C(n13762), .Y(n13759) );
  AOI22X1 U12275 ( .A(\regX[13][4] ), .B(n13259), .C(\regX[17][4] ), .D(n12803), .Y(n13762) );
  INVX1 U12276 ( .A(Out_direction[4]), .Y(n13739) );
  INVX1 U12277 ( .A(Out_gf[4]), .Y(n12527) );
  OAI21X1 U12278 ( .A(n12525), .B(n13654), .C(n13763), .Y(n4571) );
  MUX2X1 U12279 ( .B(n13764), .A(N4480), .S(n13657), .Y(n13763) );
  OAI21X1 U12280 ( .A(n13658), .B(n13765), .C(n13766), .Y(n13764) );
  AOI22X1 U12281 ( .A(n13661), .B(n13767), .C(Out_gradient[3]), .D(n13663), 
        .Y(n13766) );
  NAND3X1 U12282 ( .A(n13768), .B(n13769), .C(n13770), .Y(n13767) );
  NOR2X1 U12283 ( .A(n13771), .B(n13772), .Y(n13770) );
  OR2X1 U12284 ( .A(n13773), .B(n13774), .Y(n13772) );
  OAI21X1 U12285 ( .A(n13256), .B(n12846), .C(n13775), .Y(n13774) );
  AOI22X1 U12286 ( .A(N1378), .B(n12710), .C(\regX[19][3] ), .D(n13185), .Y(
        n13775) );
  OAI21X1 U12287 ( .A(n12723), .B(n12716), .C(n13776), .Y(n13773) );
  AOI22X1 U12288 ( .A(\regX[5][3] ), .B(n12745), .C(\regX[0][3] ), .D(n12607), 
        .Y(n13776) );
  NAND3X1 U12289 ( .A(n13777), .B(n13778), .C(n13779), .Y(n13771) );
  AOI21X1 U12290 ( .A(\regX[1][3] ), .B(n12699), .C(n13780), .Y(n13779) );
  OAI22X1 U12291 ( .A(n13271), .B(n13170), .C(n13268), .D(n12895), .Y(n13780)
         );
  AOI22X1 U12292 ( .A(\regX[9][3] ), .B(n12781), .C(\regX[8][3] ), .D(n12769), 
        .Y(n13778) );
  AOI22X1 U12293 ( .A(N1618), .B(n12890), .C(N1680), .D(n12632), .Y(n13777) );
  NOR2X1 U12294 ( .A(n13781), .B(n13782), .Y(n13769) );
  OAI21X1 U12295 ( .A(n12735), .B(n12728), .C(n13783), .Y(n13782) );
  AOI22X1 U12296 ( .A(\regX[20][3] ), .B(n12870), .C(\regX[24][3] ), .D(n12817), .Y(n13783) );
  OAI21X1 U12297 ( .A(n13253), .B(n12836), .C(n13784), .Y(n13781) );
  AOI22X1 U12298 ( .A(\regX[7][3] ), .B(n12756), .C(\regX[16][3] ), .D(n12791), 
        .Y(n13784) );
  NOR2X1 U12299 ( .A(n13785), .B(n13786), .Y(n13768) );
  OAI21X1 U12300 ( .A(n12678), .B(n12673), .C(n13787), .Y(n13786) );
  AOI22X1 U12301 ( .A(\regX[15][3] ), .B(n13250), .C(\regX[21][3] ), .D(n12880), .Y(n13787) );
  OAI21X1 U12302 ( .A(n13247), .B(n12825), .C(n13788), .Y(n13785) );
  AOI22X1 U12303 ( .A(\regX[13][3] ), .B(n13259), .C(\regX[17][3] ), .D(n12803), .Y(n13788) );
  INVX1 U12304 ( .A(Out_direction[3]), .Y(n13765) );
  INVX1 U12305 ( .A(Out_gf[3]), .Y(n12525) );
  OAI21X1 U12306 ( .A(n12523), .B(n13654), .C(n13789), .Y(n4569) );
  MUX2X1 U12307 ( .B(n13790), .A(N4483), .S(n13657), .Y(n13789) );
  OAI21X1 U12308 ( .A(n13658), .B(n13791), .C(n13792), .Y(n13790) );
  AOI22X1 U12309 ( .A(n13661), .B(n13793), .C(Out_gradient[2]), .D(n13663), 
        .Y(n13792) );
  NAND3X1 U12310 ( .A(n13794), .B(n13795), .C(n13796), .Y(n13793) );
  NOR2X1 U12311 ( .A(n13797), .B(n13798), .Y(n13796) );
  OR2X1 U12312 ( .A(n13799), .B(n13800), .Y(n13798) );
  OAI21X1 U12313 ( .A(n13256), .B(n12845), .C(n13801), .Y(n13800) );
  AOI22X1 U12314 ( .A(N1377), .B(n12710), .C(\regX[19][2] ), .D(n13185), .Y(
        n13801) );
  OAI21X1 U12315 ( .A(n12723), .B(n12715), .C(n13802), .Y(n13799) );
  AOI22X1 U12316 ( .A(\regX[5][2] ), .B(n12745), .C(\regX[0][2] ), .D(n12607), 
        .Y(n13802) );
  NAND3X1 U12317 ( .A(n13803), .B(n13804), .C(n13805), .Y(n13797) );
  AOI21X1 U12318 ( .A(\regX[1][2] ), .B(n12699), .C(n13806), .Y(n13805) );
  OAI22X1 U12319 ( .A(n13271), .B(n13169), .C(n13268), .D(n12894), .Y(n13806)
         );
  AOI22X1 U12320 ( .A(\regX[9][2] ), .B(n12781), .C(\regX[8][2] ), .D(n12769), 
        .Y(n13804) );
  AOI22X1 U12321 ( .A(N1617), .B(n12890), .C(N1679), .D(n12632), .Y(n13803) );
  NOR2X1 U12322 ( .A(n13807), .B(n13808), .Y(n13795) );
  OAI21X1 U12323 ( .A(n12735), .B(n12727), .C(n13809), .Y(n13808) );
  AOI22X1 U12324 ( .A(\regX[20][2] ), .B(n12870), .C(\regX[24][2] ), .D(n12817), .Y(n13809) );
  OAI21X1 U12325 ( .A(n13253), .B(n12835), .C(n13810), .Y(n13807) );
  AOI22X1 U12326 ( .A(\regX[7][2] ), .B(n12756), .C(\regX[16][2] ), .D(n12791), 
        .Y(n13810) );
  NOR2X1 U12327 ( .A(n13811), .B(n13812), .Y(n13794) );
  OAI21X1 U12328 ( .A(n12678), .B(n12672), .C(n13813), .Y(n13812) );
  AOI22X1 U12329 ( .A(\regX[15][2] ), .B(n13250), .C(\regX[21][2] ), .D(n12880), .Y(n13813) );
  OAI21X1 U12330 ( .A(n13247), .B(n12824), .C(n13814), .Y(n13811) );
  AOI22X1 U12331 ( .A(\regX[13][2] ), .B(n13259), .C(\regX[17][2] ), .D(n12803), .Y(n13814) );
  INVX1 U12332 ( .A(Out_direction[2]), .Y(n13791) );
  INVX1 U12333 ( .A(Out_gf[2]), .Y(n12523) );
  OAI21X1 U12334 ( .A(n12521), .B(n13654), .C(n13815), .Y(n4567) );
  MUX2X1 U12335 ( .B(n13816), .A(N4486), .S(n13657), .Y(n13815) );
  OAI21X1 U12336 ( .A(n13658), .B(n13817), .C(n13818), .Y(n13816) );
  AOI22X1 U12337 ( .A(n13661), .B(n13819), .C(Out_gradient[1]), .D(n13663), 
        .Y(n13818) );
  NAND3X1 U12338 ( .A(n13820), .B(n13821), .C(n13822), .Y(n13819) );
  NOR2X1 U12339 ( .A(n13823), .B(n13824), .Y(n13822) );
  OR2X1 U12340 ( .A(n13825), .B(n13826), .Y(n13824) );
  OAI21X1 U12341 ( .A(n13256), .B(n12844), .C(n13827), .Y(n13826) );
  AOI22X1 U12342 ( .A(N1376), .B(n12710), .C(\regX[19][1] ), .D(n13185), .Y(
        n13827) );
  OAI21X1 U12343 ( .A(n12723), .B(n12714), .C(n13828), .Y(n13825) );
  AOI22X1 U12344 ( .A(\regX[5][1] ), .B(n12745), .C(\regX[0][1] ), .D(n12607), 
        .Y(n13828) );
  NAND3X1 U12345 ( .A(n13829), .B(n13830), .C(n13831), .Y(n13823) );
  AOI21X1 U12346 ( .A(\regX[1][1] ), .B(n12699), .C(n13832), .Y(n13831) );
  OAI22X1 U12347 ( .A(n13271), .B(n13168), .C(n13268), .D(n12893), .Y(n13832)
         );
  AOI22X1 U12348 ( .A(\regX[9][1] ), .B(n12781), .C(\regX[8][1] ), .D(n12769), 
        .Y(n13830) );
  AOI22X1 U12349 ( .A(N1616), .B(n12890), .C(N1678), .D(n12632), .Y(n13829) );
  INVX1 U12350 ( .A(n13833), .Y(n12632) );
  INVX1 U12351 ( .A(n13834), .Y(n12890) );
  NOR2X1 U12352 ( .A(n13835), .B(n13836), .Y(n13821) );
  OAI21X1 U12353 ( .A(n12735), .B(n12726), .C(n13837), .Y(n13836) );
  AOI22X1 U12354 ( .A(\regX[20][1] ), .B(n12870), .C(\regX[24][1] ), .D(n12817), .Y(n13837) );
  OAI21X1 U12355 ( .A(n13253), .B(n12834), .C(n13838), .Y(n13835) );
  AOI22X1 U12356 ( .A(\regX[7][1] ), .B(n12756), .C(\regX[16][1] ), .D(n12791), 
        .Y(n13838) );
  NOR2X1 U12357 ( .A(n13839), .B(n13840), .Y(n13820) );
  OAI21X1 U12358 ( .A(n12678), .B(n12671), .C(n13841), .Y(n13840) );
  AOI22X1 U12359 ( .A(\regX[15][1] ), .B(n13250), .C(\regX[21][1] ), .D(n12880), .Y(n13841) );
  OAI21X1 U12360 ( .A(n13247), .B(n12823), .C(n13842), .Y(n13839) );
  AOI22X1 U12361 ( .A(\regX[13][1] ), .B(n13259), .C(\regX[17][1] ), .D(n12803), .Y(n13842) );
  INVX1 U12362 ( .A(Out_direction[1]), .Y(n13817) );
  INVX1 U12363 ( .A(Out_gf[1]), .Y(n12521) );
  OAI21X1 U12364 ( .A(n12518), .B(n13654), .C(n13843), .Y(n4565) );
  MUX2X1 U12365 ( .B(n13844), .A(N4489), .S(n13657), .Y(n13843) );
  NAND3X1 U12366 ( .A(n13845), .B(n13846), .C(n13847), .Y(n13844) );
  AOI22X1 U12367 ( .A(Out_gradient[0]), .B(n13663), .C(Out_direction[0]), .D(
        n13848), .Y(n13847) );
  INVX1 U12368 ( .A(n13658), .Y(n13848) );
  NAND3X1 U12369 ( .A(n12561), .B(n12564), .C(dReadReg[1]), .Y(n13658) );
  INVX1 U12370 ( .A(n13849), .Y(n13663) );
  NAND3X1 U12371 ( .A(n12561), .B(n12562), .C(dReadReg[0]), .Y(n13849) );
  INVX1 U12372 ( .A(dReadReg[1]), .Y(n12562) );
  NAND3X1 U12373 ( .A(n13850), .B(n12564), .C(n13851), .Y(n13846) );
  AND2X1 U12374 ( .A(\Out_bThres[0] ), .B(dReadReg[2]), .Y(n13851) );
  INVX1 U12375 ( .A(dReadReg[0]), .Y(n12564) );
  NOR2X1 U12376 ( .A(dReadReg[3]), .B(dReadReg[1]), .Y(n13850) );
  OAI21X1 U12377 ( .A(n13852), .B(n13853), .C(n13661), .Y(n13845) );
  INVX1 U12378 ( .A(n13854), .Y(n13661) );
  NAND3X1 U12379 ( .A(dReadReg[0]), .B(n12561), .C(dReadReg[1]), .Y(n13854) );
  NAND2X1 U12380 ( .A(n13855), .B(n13856), .Y(n13853) );
  NOR2X1 U12381 ( .A(n13857), .B(n13858), .Y(n13856) );
  OAI21X1 U12382 ( .A(n12735), .B(n12724), .C(n13859), .Y(n13858) );
  AOI22X1 U12383 ( .A(\regX[20][0] ), .B(n12870), .C(\regX[24][0] ), .D(n12817), .Y(n13859) );
  NOR2X1 U12384 ( .A(n12902), .B(n13189), .Y(n12817) );
  AND2X1 U12385 ( .A(n13860), .B(n13861), .Y(n12870) );
  NAND2X1 U12386 ( .A(n13861), .B(n13862), .Y(n12735) );
  OAI21X1 U12387 ( .A(n13253), .B(n12832), .C(n13863), .Y(n13857) );
  AOI22X1 U12388 ( .A(\regX[7][0] ), .B(n12756), .C(\regX[16][0] ), .D(n12791), 
        .Y(n13863) );
  INVX1 U12389 ( .A(n13238), .Y(n12791) );
  NAND3X1 U12390 ( .A(n12816), .B(n13189), .C(N981), .Y(n13238) );
  INVX1 U12391 ( .A(n13230), .Y(n12756) );
  NAND2X1 U12392 ( .A(n13864), .B(n13865), .Y(n13230) );
  NAND2X1 U12393 ( .A(n13860), .B(n13865), .Y(n13253) );
  NOR2X1 U12394 ( .A(n13866), .B(n13867), .Y(n13855) );
  OAI21X1 U12395 ( .A(n12678), .B(n12669), .C(n13868), .Y(n13867) );
  AOI22X1 U12396 ( .A(\regX[15][0] ), .B(n13250), .C(\regX[21][0] ), .D(n12880), .Y(n13868) );
  AND2X1 U12397 ( .A(n13869), .B(n13861), .Y(n12880) );
  INVX1 U12398 ( .A(n12594), .Y(n13250) );
  NAND2X1 U12399 ( .A(n13870), .B(n13865), .Y(n12594) );
  OAI21X1 U12400 ( .A(n13247), .B(n12821), .C(n13871), .Y(n13866) );
  AOI22X1 U12401 ( .A(\regX[13][0] ), .B(n13259), .C(\regX[17][0] ), .D(n12803), .Y(n13871) );
  NOR2X1 U12402 ( .A(n12902), .B(n13872), .Y(n12803) );
  INVX1 U12403 ( .A(n12619), .Y(n13259) );
  NAND2X1 U12404 ( .A(n13861), .B(n13870), .Y(n12619) );
  NAND2X1 U12405 ( .A(n13873), .B(n13865), .Y(n13247) );
  NAND3X1 U12406 ( .A(n13874), .B(n13875), .C(n13876), .Y(n13852) );
  NOR2X1 U12407 ( .A(n13877), .B(n13878), .Y(n13876) );
  OAI21X1 U12408 ( .A(n13256), .B(n12842), .C(n13879), .Y(n13878) );
  AOI22X1 U12409 ( .A(N1375), .B(n12710), .C(\regX[19][0] ), .D(n13185), .Y(
        n13879) );
  AND2X1 U12410 ( .A(n13869), .B(n13880), .Y(n13185) );
  INVX1 U12411 ( .A(n13276), .Y(n12710) );
  NAND2X1 U12412 ( .A(n13880), .B(n13862), .Y(n13276) );
  NAND2X1 U12413 ( .A(n13869), .B(n13865), .Y(n13256) );
  NOR2X1 U12414 ( .A(n12902), .B(n13881), .Y(n13869) );
  OAI21X1 U12415 ( .A(n12723), .B(n12712), .C(n13882), .Y(n13877) );
  AOI22X1 U12416 ( .A(\regX[5][0] ), .B(n12745), .C(\regX[0][0] ), .D(n12607), 
        .Y(n13882) );
  NOR2X1 U12417 ( .A(n13883), .B(n13884), .Y(n12607) );
  INVX1 U12418 ( .A(n13225), .Y(n12745) );
  NAND2X1 U12419 ( .A(n13864), .B(n13861), .Y(n13225) );
  NAND2X1 U12420 ( .A(n13864), .B(n13880), .Y(n12723) );
  NOR2X1 U12421 ( .A(n13881), .B(n13884), .Y(n13864) );
  NOR2X1 U12422 ( .A(n13885), .B(n13886), .Y(n13875) );
  OAI22X1 U12423 ( .A(n13833), .B(n12852), .C(n13834), .D(n12881), .Y(n13886)
         );
  NAND2X1 U12424 ( .A(n13880), .B(n13873), .Y(n13834) );
  NAND2X1 U12425 ( .A(n13873), .B(n13861), .Y(n13833) );
  NOR2X1 U12426 ( .A(n13887), .B(N978), .Y(n13861) );
  NOR2X1 U12427 ( .A(n13189), .B(N977), .Y(n13873) );
  INVX1 U12428 ( .A(n13888), .Y(n13885) );
  AOI22X1 U12429 ( .A(n12769), .B(\regX[8][0] ), .C(n12781), .D(\regX[9][0] ), 
        .Y(n13888) );
  NOR2X1 U12430 ( .A(n13872), .B(n13189), .Y(n12781) );
  INVX1 U12431 ( .A(n13233), .Y(n12769) );
  NAND3X1 U12432 ( .A(N980), .B(n12902), .C(n12816), .Y(n13233) );
  INVX1 U12433 ( .A(n13883), .Y(n12816) );
  NAND3X1 U12434 ( .A(n13889), .B(n13887), .C(n13881), .Y(n13883) );
  AOI21X1 U12435 ( .A(\regX[1][0] ), .B(n12699), .C(n13890), .Y(n13874) );
  OAI22X1 U12436 ( .A(n12555), .B(n13271), .C(n13268), .D(n12891), .Y(n13890)
         );
  NAND2X1 U12437 ( .A(n13880), .B(n13870), .Y(n13268) );
  NOR2X1 U12438 ( .A(n13189), .B(n13881), .Y(n13870) );
  INVX1 U12439 ( .A(N977), .Y(n13881) );
  NAND2X1 U12440 ( .A(n13860), .B(n13880), .Y(n13271) );
  NOR2X1 U12441 ( .A(n13889), .B(N979), .Y(n13880) );
  NOR2X1 U12442 ( .A(n12902), .B(N977), .Y(n13860) );
  NOR2X1 U12443 ( .A(n13872), .B(n13884), .Y(n12699) );
  NAND3X1 U12444 ( .A(n13889), .B(n13887), .C(N977), .Y(n13872) );
  NAND3X1 U12445 ( .A(n12561), .B(n12557), .C(n13891), .Y(n13654) );
  NOR2X1 U12446 ( .A(dReadReg[1]), .B(dReadReg[0]), .Y(n13891) );
  INVX1 U12447 ( .A(n13657), .Y(n12557) );
  NAND3X1 U12448 ( .A(rst_b), .B(n12556), .C(bWE), .Y(n13657) );
  NOR2X1 U12449 ( .A(dReadReg[2]), .B(dReadReg[3]), .Y(n12561) );
  INVX1 U12450 ( .A(Out_gf[0]), .Y(n12518) );
  INVX1 U12451 ( .A(n13894), .Y(n12459) );
  MUX2X1 U12452 ( .B(N2558), .A(Gx[0]), .S(n8303), .Y(n13894) );
  INVX1 U12453 ( .A(n13895), .Y(n12458) );
  MUX2X1 U12454 ( .B(N2559), .A(Gx[1]), .S(n8303), .Y(n13895) );
  INVX1 U12455 ( .A(n13896), .Y(n12457) );
  MUX2X1 U12456 ( .B(N2560), .A(Gx[2]), .S(n8303), .Y(n13896) );
  INVX1 U12457 ( .A(n13897), .Y(n12456) );
  MUX2X1 U12458 ( .B(N2561), .A(Gx[3]), .S(n8303), .Y(n13897) );
  INVX1 U12459 ( .A(n13898), .Y(n12455) );
  MUX2X1 U12460 ( .B(N2562), .A(Gx[4]), .S(n8303), .Y(n13898) );
  INVX1 U12461 ( .A(n13899), .Y(n12454) );
  MUX2X1 U12462 ( .B(N2563), .A(Gx[5]), .S(n8303), .Y(n13899) );
  INVX1 U12463 ( .A(n13900), .Y(n12453) );
  MUX2X1 U12464 ( .B(N2564), .A(Gx[6]), .S(n8303), .Y(n13900) );
  INVX1 U12465 ( .A(n13901), .Y(n12452) );
  MUX2X1 U12466 ( .B(N2565), .A(Gx[7]), .S(n8303), .Y(n13901) );
  INVX1 U12467 ( .A(n13902), .Y(n12451) );
  MUX2X1 U12468 ( .B(N2566), .A(Gx[8]), .S(n8303), .Y(n13902) );
  INVX1 U12469 ( .A(n13903), .Y(n12450) );
  MUX2X1 U12470 ( .B(N2567), .A(Gx[9]), .S(n8303), .Y(n13903) );
  INVX1 U12471 ( .A(n13904), .Y(n12449) );
  MUX2X1 U12472 ( .B(N2568), .A(Gx[10]), .S(n8303), .Y(n13904) );
  INVX1 U12473 ( .A(n13906), .Y(n12448) );
  MUX2X1 U12474 ( .B(N4432), .A(n13907), .S(n13196), .Y(n13906) );
  AND2X1 U12475 ( .A(n13908), .B(n12668), .Y(n13196) );
  INVX1 U12476 ( .A(n12680), .Y(n12668) );
  NAND3X1 U12477 ( .A(rst_b), .B(n12513), .C(bCE), .Y(n12680) );
  INVX1 U12478 ( .A(bOPEnable), .Y(n12513) );
  AOI21X1 U12479 ( .A(n13217), .B(n13909), .C(n12570), .Y(n13908) );
  OAI21X1 U12480 ( .A(n13907), .B(n13910), .C(n13911), .Y(n13909) );
  MUX2X1 U12481 ( .B(n13216), .A(n13209), .S(n13202), .Y(n13910) );
  INVX1 U12482 ( .A(n13215), .Y(n13202) );
  INVX1 U12483 ( .A(n13912), .Y(n13209) );
  NOR2X1 U12484 ( .A(n12471), .B(n12537), .Y(n13217) );
  OAI21X1 U12485 ( .A(n13913), .B(n13912), .C(n13212), .Y(n13907) );
  NAND3X1 U12486 ( .A(n13215), .B(n13216), .C(N2874), .Y(n13212) );
  NAND2X1 U12487 ( .A(N3336), .B(N2841), .Y(n13216) );
  NOR2X1 U12488 ( .A(n13165), .B(N2777), .Y(n13215) );
  NAND2X1 U12489 ( .A(n13165), .B(N2880), .Y(n13912) );
  NOR2X1 U12490 ( .A(N2945), .B(n12687), .Y(n13913) );
  INVX1 U12491 ( .A(n13914), .Y(n12447) );
  MUX2X1 U12492 ( .B(InData[2]), .A(\regY[6][2] ), .S(n12491), .Y(n13914) );
  INVX1 U12493 ( .A(n13915), .Y(n12446) );
  MUX2X1 U12494 ( .B(InData[0]), .A(\regY[6][0] ), .S(n12491), .Y(n13915) );
  NAND3X1 U12495 ( .A(n13193), .B(n13192), .C(n13916), .Y(n12491) );
  NOR2X1 U12496 ( .A(n12678), .B(n13191), .Y(n13916) );
  INVX1 U12497 ( .A(dWriteReg[0]), .Y(n13191) );
  NAND2X1 U12498 ( .A(n13865), .B(n13862), .Y(n12678) );
  NOR2X1 U12499 ( .A(n13884), .B(N977), .Y(n13862) );
  NAND2X1 U12500 ( .A(n13189), .B(n12902), .Y(n13884) );
  INVX1 U12501 ( .A(N981), .Y(n12902) );
  INVX1 U12502 ( .A(N980), .Y(n13189) );
  NOR2X1 U12503 ( .A(n13887), .B(n13889), .Y(n13865) );
  INVX1 U12504 ( .A(N978), .Y(n13889) );
  INVX1 U12505 ( .A(N979), .Y(n13887) );
  INVX1 U12506 ( .A(dWriteReg[1]), .Y(n13192) );
  INVX1 U12507 ( .A(n13917), .Y(n13193) );
  NAND3X1 U12508 ( .A(n13283), .B(n13285), .C(rst_b), .Y(n13917) );
  NOR2X1 U12509 ( .A(dWriteReg[2]), .B(dWriteReg[3]), .Y(n13285) );
  INVX1 U12510 ( .A(n13281), .Y(n13283) );
  NAND3X1 U12511 ( .A(n13194), .B(n13195), .C(n12494), .Y(n13281) );
  NOR2X1 U12512 ( .A(bCE), .B(bWE), .Y(n12494) );
  INVX1 U12513 ( .A(N983), .Y(n13195) );
  INVX1 U12514 ( .A(N982), .Y(n13194) );
  OAI21X1 U12515 ( .A(n12470), .B(n12879), .C(n13918), .Y(\U3/U98/Z_7 ) );
  OAI21X1 U12516 ( .A(n12470), .B(n12878), .C(n13918), .Y(\U3/U98/Z_6 ) );
  OAI21X1 U12517 ( .A(n12470), .B(n12877), .C(n13918), .Y(\U3/U98/Z_5 ) );
  OAI21X1 U12518 ( .A(n12470), .B(n12876), .C(n13918), .Y(\U3/U98/Z_4 ) );
  OAI21X1 U12519 ( .A(n12470), .B(n12875), .C(n13918), .Y(\U3/U98/Z_3 ) );
  OAI21X1 U12520 ( .A(n12470), .B(n12874), .C(n13918), .Y(\U3/U98/Z_2 ) );
  OAI21X1 U12521 ( .A(n12470), .B(n12873), .C(n13918), .Y(\U3/U98/Z_1 ) );
  NAND2X1 U12522 ( .A(dy[1]), .B(n15327), .Y(n13918) );
  OAI22X1 U12523 ( .A(n12553), .B(n13405), .C(n12470), .D(n12871), .Y(
        \U3/U98/Z_0 ) );
  NAND2X1 U12524 ( .A(n13405), .B(n12470), .Y(\U3/U97/Z_0 ) );
  NAND2X1 U12525 ( .A(n12474), .B(n12464), .Y(\U3/U96/Z_0 ) );
  NAND2X1 U12526 ( .A(n13921), .B(n12464), .Y(\U3/U95/Z_0 ) );
  AND2X1 U12527 ( .A(N2890), .B(n12466), .Y(\U3/U94/Z_9 ) );
  AND2X1 U12528 ( .A(N2889), .B(n12466), .Y(\U3/U94/Z_8 ) );
  OAI21X1 U12529 ( .A(n13921), .B(n12677), .C(n13922), .Y(\U3/U94/Z_7 ) );
  NAND2X1 U12530 ( .A(N2888), .B(n12466), .Y(n13922) );
  OAI21X1 U12531 ( .A(n13921), .B(n12676), .C(n13923), .Y(\U3/U94/Z_6 ) );
  NAND2X1 U12532 ( .A(N2887), .B(n12466), .Y(n13923) );
  OAI21X1 U12533 ( .A(n13921), .B(n12675), .C(n13924), .Y(\U3/U94/Z_5 ) );
  NAND2X1 U12534 ( .A(N2886), .B(n12466), .Y(n13924) );
  OAI21X1 U12535 ( .A(n13921), .B(n12674), .C(n13925), .Y(\U3/U94/Z_4 ) );
  NAND2X1 U12536 ( .A(N2885), .B(n12466), .Y(n13925) );
  NOR2X1 U12537 ( .A(n12464), .B(n13926), .Y(\U3/U94/Z_31 ) );
  OAI21X1 U12538 ( .A(n12673), .B(n13921), .C(n13927), .Y(\U3/U94/Z_3 ) );
  NAND2X1 U12539 ( .A(N2884), .B(n12466), .Y(n13927) );
  NOR2X1 U12540 ( .A(n12464), .B(n13928), .Y(\U3/U94/Z_29 ) );
  NOR2X1 U12541 ( .A(n12464), .B(n13929), .Y(\U3/U94/Z_28 ) );
  NOR2X1 U12542 ( .A(n12464), .B(n13930), .Y(\U3/U94/Z_27 ) );
  NOR2X1 U12543 ( .A(n12464), .B(n13931), .Y(\U3/U94/Z_26 ) );
  NOR2X1 U12544 ( .A(n12464), .B(n13932), .Y(\U3/U94/Z_25 ) );
  NOR2X1 U12545 ( .A(n12464), .B(n13933), .Y(\U3/U94/Z_24 ) );
  NOR2X1 U12546 ( .A(n12464), .B(n13934), .Y(\U3/U94/Z_23 ) );
  NOR2X1 U12547 ( .A(n12464), .B(n13935), .Y(\U3/U94/Z_22 ) );
  NOR2X1 U12548 ( .A(n12464), .B(n13936), .Y(\U3/U94/Z_21 ) );
  NOR2X1 U12549 ( .A(n12464), .B(n13937), .Y(\U3/U94/Z_20 ) );
  OAI21X1 U12550 ( .A(n12672), .B(n13921), .C(n13938), .Y(\U3/U94/Z_2 ) );
  NAND2X1 U12551 ( .A(N2883), .B(n12466), .Y(n13938) );
  NOR2X1 U12552 ( .A(n12464), .B(n13939), .Y(\U3/U94/Z_19 ) );
  NOR2X1 U12553 ( .A(n12464), .B(n13940), .Y(\U3/U94/Z_18 ) );
  NOR2X1 U12554 ( .A(n12464), .B(n13941), .Y(\U3/U94/Z_17 ) );
  NOR2X1 U12555 ( .A(n13920), .B(n13942), .Y(\U3/U94/Z_16 ) );
  NOR2X1 U12556 ( .A(n12464), .B(n13943), .Y(\U3/U94/Z_15 ) );
  NOR2X1 U12557 ( .A(n13920), .B(n13944), .Y(\U3/U94/Z_14 ) );
  AND2X1 U12558 ( .A(N2894), .B(n12466), .Y(\U3/U94/Z_13 ) );
  AND2X1 U12559 ( .A(N2893), .B(n12466), .Y(\U3/U94/Z_12 ) );
  AND2X1 U12560 ( .A(N2892), .B(n12466), .Y(\U3/U94/Z_11 ) );
  AND2X1 U12561 ( .A(N2891), .B(n12466), .Y(\U3/U94/Z_10 ) );
  OAI21X1 U12562 ( .A(n12671), .B(n13921), .C(n13945), .Y(\U3/U94/Z_1 ) );
  NAND2X1 U12563 ( .A(N2882), .B(n12466), .Y(n13945) );
  OAI21X1 U12564 ( .A(n12669), .B(n13921), .C(n13946), .Y(\U3/U94/Z_0 ) );
  NAND2X1 U12565 ( .A(N2881), .B(n12466), .Y(n13946) );
  OAI21X1 U12566 ( .A(n13061), .B(n12474), .C(n13947), .Y(\U3/U93/Z_9 ) );
  INVX1 U12567 ( .A(n15332), .Y(n13947) );
  NOR2X1 U12568 ( .A(n12986), .B(n12464), .Y(n15332) );
  OAI21X1 U12569 ( .A(n13059), .B(n12474), .C(n13948), .Y(\U3/U93/Z_8 ) );
  INVX1 U12570 ( .A(n15333), .Y(n13948) );
  NOR2X1 U12571 ( .A(n12984), .B(n13920), .Y(n15333) );
  OAI21X1 U12572 ( .A(n13055), .B(n12474), .C(n13949), .Y(\U3/U93/Z_7 ) );
  AOI21X1 U12573 ( .A(n15369), .B(n13950), .C(\U3/U121/Z_7 ), .Y(n13949) );
  NAND3X1 U12574 ( .A(n13951), .B(n13952), .C(n13953), .Y(n13950) );
  NOR2X1 U12575 ( .A(n13954), .B(n13955), .Y(n13953) );
  OR2X1 U12576 ( .A(n13956), .B(n13957), .Y(n13955) );
  OAI21X1 U12577 ( .A(n12860), .B(n13958), .C(n13959), .Y(n13957) );
  AOI22X1 U12578 ( .A(n13960), .B(\regX[16][7] ), .C(n13961), .D(\regX[20][7] ), .Y(n13959) );
  OAI21X1 U12579 ( .A(n12610), .B(n13962), .C(n13963), .Y(n13956) );
  AOI22X1 U12580 ( .A(n13964), .B(N1742), .C(n13965), .D(\regX[19][7] ), .Y(
        n13963) );
  INVX1 U12581 ( .A(\regX[13][7] ), .Y(n12610) );
  NAND3X1 U12582 ( .A(n13966), .B(n13967), .C(n13968), .Y(n13954) );
  AOI21X1 U12583 ( .A(n13969), .B(\regX[15][7] ), .C(n13970), .Y(n13968) );
  OAI22X1 U12584 ( .A(n12812), .B(n13971), .C(n12850), .D(n13972), .Y(n13970)
         );
  AOI22X1 U12585 ( .A(n13973), .B(\regX[18][7] ), .C(n13974), .D(\regX[21][7] ), .Y(n13967) );
  AOI22X1 U12586 ( .A(n13975), .B(\regX[22][7] ), .C(n13976), .D(\regX[17][7] ), .Y(n13966) );
  NOR2X1 U12587 ( .A(n13977), .B(n13978), .Y(n13952) );
  OAI21X1 U12588 ( .A(n12677), .B(n13979), .C(n13980), .Y(n13978) );
  AOI22X1 U12589 ( .A(n13981), .B(\regX[8][7] ), .C(n13982), .D(\regX[7][7] ), 
        .Y(n13980) );
  OAI21X1 U12590 ( .A(n12779), .B(n13983), .C(n13984), .Y(n13977) );
  AOI22X1 U12591 ( .A(n13985), .B(\regX[11][7] ), .C(n13986), .D(N1622), .Y(
        n13984) );
  NOR2X1 U12592 ( .A(n13987), .B(n13988), .Y(n13951) );
  OAI21X1 U12593 ( .A(n12603), .B(n13989), .C(n13990), .Y(n13988) );
  AOI22X1 U12594 ( .A(n13991), .B(N1382), .C(n13992), .D(\regX[1][7] ), .Y(
        n13990) );
  OAI21X1 U12595 ( .A(n12720), .B(n13993), .C(n13994), .Y(n13987) );
  AOI22X1 U12596 ( .A(n13995), .B(\regX[5][7] ), .C(n13996), .D(N1440), .Y(
        n13994) );
  OAI21X1 U12597 ( .A(n13052), .B(n12474), .C(n13997), .Y(\U3/U93/Z_6 ) );
  AOI21X1 U12598 ( .A(n15369), .B(n13998), .C(\U3/U121/Z_6 ), .Y(n13997) );
  NAND3X1 U12599 ( .A(n13999), .B(n14000), .C(n14001), .Y(n13998) );
  NOR2X1 U12600 ( .A(n14002), .B(n14003), .Y(n14001) );
  OR2X1 U12601 ( .A(n14004), .B(n14005), .Y(n14003) );
  OAI21X1 U12602 ( .A(n12859), .B(n13958), .C(n14006), .Y(n14005) );
  AOI22X1 U12603 ( .A(n13960), .B(\regX[16][6] ), .C(n13961), .D(\regX[20][6] ), .Y(n14006) );
  OAI21X1 U12604 ( .A(n12612), .B(n13962), .C(n14007), .Y(n14004) );
  AOI22X1 U12605 ( .A(n13964), .B(N1741), .C(n13965), .D(\regX[19][6] ), .Y(
        n14007) );
  INVX1 U12606 ( .A(\regX[13][6] ), .Y(n12612) );
  NAND3X1 U12607 ( .A(n14008), .B(n14009), .C(n14010), .Y(n14002) );
  AOI21X1 U12608 ( .A(n13969), .B(\regX[15][6] ), .C(n14011), .Y(n14010) );
  OAI22X1 U12609 ( .A(n12811), .B(n13971), .C(n12849), .D(n13972), .Y(n14011)
         );
  AOI22X1 U12610 ( .A(n13973), .B(\regX[18][6] ), .C(n13974), .D(\regX[21][6] ), .Y(n14009) );
  AOI22X1 U12611 ( .A(n13975), .B(\regX[22][6] ), .C(n13976), .D(\regX[17][6] ), .Y(n14008) );
  NOR2X1 U12612 ( .A(n14012), .B(n14013), .Y(n14000) );
  OAI21X1 U12613 ( .A(n12676), .B(n13979), .C(n14014), .Y(n14013) );
  AOI22X1 U12614 ( .A(n13981), .B(\regX[8][6] ), .C(n13982), .D(\regX[7][6] ), 
        .Y(n14014) );
  OAI21X1 U12615 ( .A(n12778), .B(n13983), .C(n14015), .Y(n14012) );
  AOI22X1 U12616 ( .A(n13985), .B(\regX[11][6] ), .C(n13986), .D(N1621), .Y(
        n14015) );
  NOR2X1 U12617 ( .A(n14016), .B(n14017), .Y(n13999) );
  OAI21X1 U12618 ( .A(n12602), .B(n13989), .C(n14018), .Y(n14017) );
  AOI22X1 U12619 ( .A(n13991), .B(N1381), .C(n13992), .D(\regX[1][6] ), .Y(
        n14018) );
  OAI21X1 U12620 ( .A(n12719), .B(n13993), .C(n14019), .Y(n14016) );
  AOI22X1 U12621 ( .A(n13995), .B(\regX[5][6] ), .C(n13996), .D(N1439), .Y(
        n14019) );
  OAI21X1 U12622 ( .A(n13049), .B(n12474), .C(n14020), .Y(\U3/U93/Z_5 ) );
  AOI21X1 U12623 ( .A(n15369), .B(n14021), .C(\U3/U121/Z_5 ), .Y(n14020) );
  NAND3X1 U12624 ( .A(n14022), .B(n14023), .C(n14024), .Y(n14021) );
  NOR2X1 U12625 ( .A(n14025), .B(n14026), .Y(n14024) );
  OR2X1 U12626 ( .A(n14027), .B(n14028), .Y(n14026) );
  OAI21X1 U12627 ( .A(n12858), .B(n13958), .C(n14029), .Y(n14028) );
  AOI22X1 U12628 ( .A(n13960), .B(\regX[16][5] ), .C(n13961), .D(\regX[20][5] ), .Y(n14029) );
  OAI21X1 U12629 ( .A(n12613), .B(n13962), .C(n14030), .Y(n14027) );
  AOI22X1 U12630 ( .A(n13964), .B(N1740), .C(n13965), .D(\regX[19][5] ), .Y(
        n14030) );
  INVX1 U12631 ( .A(\regX[13][5] ), .Y(n12613) );
  NAND3X1 U12632 ( .A(n14031), .B(n14032), .C(n14033), .Y(n14025) );
  AOI21X1 U12633 ( .A(n13969), .B(\regX[15][5] ), .C(n14034), .Y(n14033) );
  OAI22X1 U12634 ( .A(n12810), .B(n13971), .C(n12848), .D(n13972), .Y(n14034)
         );
  AOI22X1 U12635 ( .A(n13973), .B(\regX[18][5] ), .C(n13974), .D(\regX[21][5] ), .Y(n14032) );
  AOI22X1 U12636 ( .A(n13975), .B(\regX[22][5] ), .C(n13976), .D(\regX[17][5] ), .Y(n14031) );
  NOR2X1 U12637 ( .A(n14035), .B(n14036), .Y(n14023) );
  OAI21X1 U12638 ( .A(n12675), .B(n13979), .C(n14037), .Y(n14036) );
  AOI22X1 U12639 ( .A(n13981), .B(\regX[8][5] ), .C(n13982), .D(\regX[7][5] ), 
        .Y(n14037) );
  OAI21X1 U12640 ( .A(n12777), .B(n13983), .C(n14038), .Y(n14035) );
  AOI22X1 U12641 ( .A(n13985), .B(\regX[11][5] ), .C(n13986), .D(N1620), .Y(
        n14038) );
  NOR2X1 U12642 ( .A(n14039), .B(n14040), .Y(n14022) );
  OAI21X1 U12643 ( .A(n12601), .B(n13989), .C(n14041), .Y(n14040) );
  AOI22X1 U12644 ( .A(n13991), .B(N1380), .C(n13992), .D(\regX[1][5] ), .Y(
        n14041) );
  OAI21X1 U12645 ( .A(n12718), .B(n13993), .C(n14042), .Y(n14039) );
  AOI22X1 U12646 ( .A(n13995), .B(\regX[5][5] ), .C(n13996), .D(N1438), .Y(
        n14042) );
  OAI21X1 U12647 ( .A(n13046), .B(n12474), .C(n14043), .Y(\U3/U93/Z_4 ) );
  AOI21X1 U12648 ( .A(n15369), .B(n14044), .C(\U3/U121/Z_4 ), .Y(n14043) );
  NAND3X1 U12649 ( .A(n14045), .B(n14046), .C(n14047), .Y(n14044) );
  NOR2X1 U12650 ( .A(n14048), .B(n14049), .Y(n14047) );
  OR2X1 U12651 ( .A(n14050), .B(n14051), .Y(n14049) );
  OAI21X1 U12652 ( .A(n12857), .B(n13958), .C(n14052), .Y(n14051) );
  AOI22X1 U12653 ( .A(n13960), .B(\regX[16][4] ), .C(n13961), .D(\regX[20][4] ), .Y(n14052) );
  OAI21X1 U12654 ( .A(n12614), .B(n13962), .C(n14053), .Y(n14050) );
  AOI22X1 U12655 ( .A(n13964), .B(N1739), .C(n13965), .D(\regX[19][4] ), .Y(
        n14053) );
  INVX1 U12656 ( .A(\regX[13][4] ), .Y(n12614) );
  NAND3X1 U12657 ( .A(n14054), .B(n14055), .C(n14056), .Y(n14048) );
  AOI21X1 U12658 ( .A(n13969), .B(\regX[15][4] ), .C(n14057), .Y(n14056) );
  OAI22X1 U12659 ( .A(n12809), .B(n13971), .C(n12847), .D(n13972), .Y(n14057)
         );
  AOI22X1 U12660 ( .A(n13973), .B(\regX[18][4] ), .C(n13974), .D(\regX[21][4] ), .Y(n14055) );
  AOI22X1 U12661 ( .A(n13975), .B(\regX[22][4] ), .C(n13976), .D(\regX[17][4] ), .Y(n14054) );
  NOR2X1 U12662 ( .A(n14058), .B(n14059), .Y(n14046) );
  OAI21X1 U12663 ( .A(n12674), .B(n13979), .C(n14060), .Y(n14059) );
  AOI22X1 U12664 ( .A(n13981), .B(\regX[8][4] ), .C(n13982), .D(\regX[7][4] ), 
        .Y(n14060) );
  OAI21X1 U12665 ( .A(n12776), .B(n13983), .C(n14061), .Y(n14058) );
  AOI22X1 U12666 ( .A(n13985), .B(\regX[11][4] ), .C(n13986), .D(N1619), .Y(
        n14061) );
  NOR2X1 U12667 ( .A(n14062), .B(n14063), .Y(n14045) );
  OAI21X1 U12668 ( .A(n12600), .B(n13989), .C(n14064), .Y(n14063) );
  AOI22X1 U12669 ( .A(n13991), .B(N1379), .C(n13992), .D(\regX[1][4] ), .Y(
        n14064) );
  OAI21X1 U12670 ( .A(n12717), .B(n13993), .C(n14065), .Y(n14062) );
  AOI22X1 U12671 ( .A(n13995), .B(\regX[5][4] ), .C(n13996), .D(N1437), .Y(
        n14065) );
  OAI21X1 U12672 ( .A(n13161), .B(n12474), .C(n14066), .Y(\U3/U93/Z_31 ) );
  INVX1 U12673 ( .A(n15334), .Y(n14066) );
  NOR2X1 U12674 ( .A(n13030), .B(n12464), .Y(n15334) );
  OAI21X1 U12675 ( .A(n13157), .B(n12474), .C(n14067), .Y(\U3/U93/Z_30 ) );
  INVX1 U12676 ( .A(n15335), .Y(n14067) );
  NOR2X1 U12677 ( .A(n13028), .B(n13920), .Y(n15335) );
  OAI21X1 U12678 ( .A(n13043), .B(n12474), .C(n14068), .Y(\U3/U93/Z_3 ) );
  AOI22X1 U12679 ( .A(n15369), .B(n14069), .C(fGy[3]), .D(n12466), .Y(n14068)
         );
  NAND3X1 U12680 ( .A(n14070), .B(n14071), .C(n14072), .Y(n14069) );
  NOR2X1 U12681 ( .A(n14073), .B(n14074), .Y(n14072) );
  OR2X1 U12682 ( .A(n14075), .B(n14076), .Y(n14074) );
  OAI21X1 U12683 ( .A(n12856), .B(n13958), .C(n14077), .Y(n14076) );
  AOI22X1 U12684 ( .A(n13960), .B(\regX[16][3] ), .C(n13961), .D(\regX[20][3] ), .Y(n14077) );
  OAI21X1 U12685 ( .A(n12615), .B(n13962), .C(n14078), .Y(n14075) );
  AOI22X1 U12686 ( .A(n13964), .B(N1738), .C(n13965), .D(\regX[19][3] ), .Y(
        n14078) );
  INVX1 U12687 ( .A(\regX[13][3] ), .Y(n12615) );
  NAND3X1 U12688 ( .A(n14079), .B(n14080), .C(n14081), .Y(n14073) );
  AOI21X1 U12689 ( .A(n13969), .B(\regX[15][3] ), .C(n14082), .Y(n14081) );
  OAI22X1 U12690 ( .A(n12808), .B(n13971), .C(n12846), .D(n13972), .Y(n14082)
         );
  AOI22X1 U12691 ( .A(n13973), .B(\regX[18][3] ), .C(n13974), .D(\regX[21][3] ), .Y(n14080) );
  AOI22X1 U12692 ( .A(n13975), .B(\regX[22][3] ), .C(n13976), .D(\regX[17][3] ), .Y(n14079) );
  NOR2X1 U12693 ( .A(n14083), .B(n14084), .Y(n14071) );
  OAI21X1 U12694 ( .A(n12673), .B(n13979), .C(n14085), .Y(n14084) );
  AOI22X1 U12695 ( .A(n13981), .B(\regX[8][3] ), .C(n13982), .D(\regX[7][3] ), 
        .Y(n14085) );
  OAI21X1 U12696 ( .A(n12775), .B(n13983), .C(n14086), .Y(n14083) );
  AOI22X1 U12697 ( .A(n13985), .B(\regX[11][3] ), .C(n13986), .D(N1618), .Y(
        n14086) );
  NOR2X1 U12698 ( .A(n14087), .B(n14088), .Y(n14070) );
  OAI21X1 U12699 ( .A(n12599), .B(n13989), .C(n14089), .Y(n14088) );
  AOI22X1 U12700 ( .A(n13991), .B(N1378), .C(n13992), .D(\regX[1][3] ), .Y(
        n14089) );
  INVX1 U12701 ( .A(\regX[0][3] ), .Y(n12599) );
  OAI21X1 U12702 ( .A(n12716), .B(n13993), .C(n14090), .Y(n14087) );
  AOI22X1 U12703 ( .A(n13995), .B(\regX[5][3] ), .C(n13996), .D(N1436), .Y(
        n14090) );
  OAI21X1 U12704 ( .A(n13153), .B(n12474), .C(n14091), .Y(\U3/U93/Z_29 ) );
  INVX1 U12705 ( .A(n15336), .Y(n14091) );
  NOR2X1 U12706 ( .A(n13026), .B(n12464), .Y(n15336) );
  OAI21X1 U12707 ( .A(n13149), .B(n12474), .C(n14092), .Y(\U3/U93/Z_28 ) );
  INVX1 U12708 ( .A(n15337), .Y(n14092) );
  NOR2X1 U12709 ( .A(n13024), .B(n13920), .Y(n15337) );
  OAI21X1 U12710 ( .A(n13145), .B(n12474), .C(n14093), .Y(\U3/U93/Z_27 ) );
  INVX1 U12711 ( .A(n15338), .Y(n14093) );
  NOR2X1 U12712 ( .A(n13022), .B(n12464), .Y(n15338) );
  OAI21X1 U12713 ( .A(n13141), .B(n12474), .C(n14094), .Y(\U3/U93/Z_26 ) );
  INVX1 U12714 ( .A(n15339), .Y(n14094) );
  NOR2X1 U12715 ( .A(n13020), .B(n13920), .Y(n15339) );
  OAI21X1 U12716 ( .A(n13137), .B(n12474), .C(n14095), .Y(\U3/U93/Z_25 ) );
  INVX1 U12717 ( .A(n15340), .Y(n14095) );
  NOR2X1 U12718 ( .A(n13018), .B(n12464), .Y(n15340) );
  OAI21X1 U12719 ( .A(n13133), .B(n12474), .C(n14096), .Y(\U3/U93/Z_24 ) );
  INVX1 U12720 ( .A(n15341), .Y(n14096) );
  NOR2X1 U12721 ( .A(n13016), .B(n13920), .Y(n15341) );
  OAI21X1 U12722 ( .A(n13129), .B(n12474), .C(n14097), .Y(\U3/U93/Z_23 ) );
  INVX1 U12723 ( .A(n15342), .Y(n14097) );
  NOR2X1 U12724 ( .A(n13014), .B(n12464), .Y(n15342) );
  OAI21X1 U12725 ( .A(n13125), .B(n12474), .C(n14098), .Y(\U3/U93/Z_22 ) );
  INVX1 U12726 ( .A(n15343), .Y(n14098) );
  NOR2X1 U12727 ( .A(n13012), .B(n13920), .Y(n15343) );
  OAI21X1 U12728 ( .A(n13121), .B(n12474), .C(n14099), .Y(\U3/U93/Z_21 ) );
  INVX1 U12729 ( .A(n15344), .Y(n14099) );
  NOR2X1 U12730 ( .A(n13010), .B(n12464), .Y(n15344) );
  OAI21X1 U12731 ( .A(n13117), .B(n12474), .C(n14100), .Y(\U3/U93/Z_20 ) );
  INVX1 U12732 ( .A(n15345), .Y(n14100) );
  NOR2X1 U12733 ( .A(n13008), .B(n13920), .Y(n15345) );
  OAI21X1 U12734 ( .A(n13040), .B(n12474), .C(n14101), .Y(\U3/U93/Z_2 ) );
  AOI22X1 U12735 ( .A(n15369), .B(n14102), .C(fGy[2]), .D(n12466), .Y(n14101)
         );
  NAND3X1 U12736 ( .A(n14103), .B(n14104), .C(n14105), .Y(n14102) );
  NOR2X1 U12737 ( .A(n14106), .B(n14107), .Y(n14105) );
  OR2X1 U12738 ( .A(n14108), .B(n14109), .Y(n14107) );
  OAI21X1 U12739 ( .A(n12855), .B(n13958), .C(n14110), .Y(n14109) );
  AOI22X1 U12740 ( .A(n13960), .B(\regX[16][2] ), .C(n13961), .D(\regX[20][2] ), .Y(n14110) );
  OAI21X1 U12741 ( .A(n12616), .B(n13962), .C(n14111), .Y(n14108) );
  AOI22X1 U12742 ( .A(n13964), .B(N1737), .C(n13965), .D(\regX[19][2] ), .Y(
        n14111) );
  INVX1 U12743 ( .A(\regX[13][2] ), .Y(n12616) );
  NAND3X1 U12744 ( .A(n14112), .B(n14113), .C(n14114), .Y(n14106) );
  AOI21X1 U12745 ( .A(n13969), .B(\regX[15][2] ), .C(n14115), .Y(n14114) );
  OAI22X1 U12746 ( .A(n12807), .B(n13971), .C(n12845), .D(n13972), .Y(n14115)
         );
  AOI22X1 U12747 ( .A(n13973), .B(\regX[18][2] ), .C(n13974), .D(\regX[21][2] ), .Y(n14113) );
  AOI22X1 U12748 ( .A(n13975), .B(\regX[22][2] ), .C(n13976), .D(\regX[17][2] ), .Y(n14112) );
  NOR2X1 U12749 ( .A(n14116), .B(n14117), .Y(n14104) );
  OAI21X1 U12750 ( .A(n12672), .B(n13979), .C(n14118), .Y(n14117) );
  AOI22X1 U12751 ( .A(n13981), .B(\regX[8][2] ), .C(n13982), .D(\regX[7][2] ), 
        .Y(n14118) );
  OAI21X1 U12752 ( .A(n12774), .B(n13983), .C(n14119), .Y(n14116) );
  AOI22X1 U12753 ( .A(n13985), .B(\regX[11][2] ), .C(n13986), .D(N1617), .Y(
        n14119) );
  NOR2X1 U12754 ( .A(n14120), .B(n14121), .Y(n14103) );
  OAI21X1 U12755 ( .A(n12597), .B(n13989), .C(n14122), .Y(n14121) );
  AOI22X1 U12756 ( .A(n13991), .B(N1377), .C(n13992), .D(\regX[1][2] ), .Y(
        n14122) );
  INVX1 U12757 ( .A(\regX[0][2] ), .Y(n12597) );
  OAI21X1 U12758 ( .A(n12715), .B(n13993), .C(n14123), .Y(n14120) );
  AOI22X1 U12759 ( .A(n13995), .B(\regX[5][2] ), .C(n13996), .D(N1435), .Y(
        n14123) );
  OAI21X1 U12760 ( .A(n13113), .B(n12474), .C(n14124), .Y(\U3/U93/Z_19 ) );
  INVX1 U12761 ( .A(n15346), .Y(n14124) );
  NOR2X1 U12762 ( .A(n13006), .B(n12464), .Y(n15346) );
  OAI21X1 U12763 ( .A(n13109), .B(n12474), .C(n14125), .Y(\U3/U93/Z_18 ) );
  INVX1 U12764 ( .A(n15347), .Y(n14125) );
  NOR2X1 U12765 ( .A(n13004), .B(n13920), .Y(n15347) );
  OAI21X1 U12766 ( .A(n13105), .B(n12474), .C(n14126), .Y(\U3/U93/Z_17 ) );
  INVX1 U12767 ( .A(n15348), .Y(n14126) );
  NOR2X1 U12768 ( .A(n13002), .B(n12464), .Y(n15348) );
  OAI21X1 U12769 ( .A(n13101), .B(n12474), .C(n14127), .Y(\U3/U93/Z_16 ) );
  INVX1 U12770 ( .A(n15349), .Y(n14127) );
  NOR2X1 U12771 ( .A(n13000), .B(n13920), .Y(n15349) );
  OAI21X1 U12772 ( .A(n13097), .B(n12474), .C(n14128), .Y(\U3/U93/Z_15 ) );
  INVX1 U12773 ( .A(n15350), .Y(n14128) );
  NOR2X1 U12774 ( .A(n12998), .B(n12464), .Y(n15350) );
  OAI21X1 U12775 ( .A(n13093), .B(n12474), .C(n14129), .Y(\U3/U93/Z_14 ) );
  INVX1 U12776 ( .A(n15351), .Y(n14129) );
  NOR2X1 U12777 ( .A(n12996), .B(n13920), .Y(n15351) );
  OAI21X1 U12778 ( .A(n13089), .B(n12474), .C(n14130), .Y(\U3/U93/Z_13 ) );
  INVX1 U12779 ( .A(n15352), .Y(n14130) );
  NOR2X1 U12780 ( .A(n12994), .B(n12464), .Y(n15352) );
  OAI21X1 U12781 ( .A(n13085), .B(n12474), .C(n14131), .Y(\U3/U93/Z_12 ) );
  INVX1 U12782 ( .A(n15353), .Y(n14131) );
  NOR2X1 U12783 ( .A(n12992), .B(n13920), .Y(n15353) );
  OAI21X1 U12784 ( .A(n13081), .B(n12474), .C(n14132), .Y(\U3/U93/Z_11 ) );
  INVX1 U12785 ( .A(n15354), .Y(n14132) );
  NOR2X1 U12786 ( .A(n12990), .B(n12464), .Y(n15354) );
  OAI21X1 U12787 ( .A(n13065), .B(n12474), .C(n14133), .Y(\U3/U93/Z_10 ) );
  INVX1 U12788 ( .A(n15355), .Y(n14133) );
  NOR2X1 U12789 ( .A(n12988), .B(n13920), .Y(n15355) );
  OAI21X1 U12790 ( .A(n13037), .B(n12474), .C(n14134), .Y(\U3/U93/Z_1 ) );
  AOI22X1 U12791 ( .A(n15369), .B(n14135), .C(fGy[1]), .D(n12466), .Y(n14134)
         );
  NAND3X1 U12792 ( .A(n14136), .B(n14137), .C(n14138), .Y(n14135) );
  NOR2X1 U12793 ( .A(n14139), .B(n14140), .Y(n14138) );
  OR2X1 U12794 ( .A(n14141), .B(n14142), .Y(n14140) );
  OAI21X1 U12795 ( .A(n12854), .B(n13958), .C(n14143), .Y(n14142) );
  AOI22X1 U12796 ( .A(n13960), .B(\regX[16][1] ), .C(n13961), .D(\regX[20][1] ), .Y(n14143) );
  OAI21X1 U12797 ( .A(n12617), .B(n13962), .C(n14144), .Y(n14141) );
  AOI22X1 U12798 ( .A(n13964), .B(N1736), .C(n13965), .D(\regX[19][1] ), .Y(
        n14144) );
  INVX1 U12799 ( .A(\regX[13][1] ), .Y(n12617) );
  NAND3X1 U12800 ( .A(n14145), .B(n14146), .C(n14147), .Y(n14139) );
  AOI21X1 U12801 ( .A(n13969), .B(\regX[15][1] ), .C(n14148), .Y(n14147) );
  OAI22X1 U12802 ( .A(n12806), .B(n13971), .C(n12844), .D(n13972), .Y(n14148)
         );
  AOI22X1 U12803 ( .A(n13973), .B(\regX[18][1] ), .C(n13974), .D(\regX[21][1] ), .Y(n14146) );
  AOI22X1 U12804 ( .A(n13975), .B(\regX[22][1] ), .C(n13976), .D(\regX[17][1] ), .Y(n14145) );
  NOR2X1 U12805 ( .A(n14149), .B(n14150), .Y(n14137) );
  OAI21X1 U12806 ( .A(n12671), .B(n13979), .C(n14151), .Y(n14150) );
  AOI22X1 U12807 ( .A(n13981), .B(\regX[8][1] ), .C(n13982), .D(\regX[7][1] ), 
        .Y(n14151) );
  OAI21X1 U12808 ( .A(n12773), .B(n13983), .C(n14152), .Y(n14149) );
  AOI22X1 U12809 ( .A(n13985), .B(\regX[11][1] ), .C(n13986), .D(N1616), .Y(
        n14152) );
  NOR2X1 U12810 ( .A(n14153), .B(n14154), .Y(n14136) );
  OAI21X1 U12811 ( .A(n12604), .B(n13989), .C(n14155), .Y(n14154) );
  AOI22X1 U12812 ( .A(n13991), .B(N1376), .C(n13992), .D(\regX[1][1] ), .Y(
        n14155) );
  INVX1 U12813 ( .A(\regX[0][1] ), .Y(n12604) );
  OAI21X1 U12814 ( .A(n12714), .B(n13993), .C(n14156), .Y(n14153) );
  AOI22X1 U12815 ( .A(n13995), .B(\regX[5][1] ), .C(n13996), .D(N1434), .Y(
        n14156) );
  OAI21X1 U12816 ( .A(n13033), .B(n12474), .C(n14157), .Y(\U3/U93/Z_0 ) );
  AOI22X1 U12817 ( .A(n15369), .B(n14158), .C(fGy[0]), .D(n12466), .Y(n14157)
         );
  NAND3X1 U12818 ( .A(n14159), .B(n14160), .C(n14161), .Y(n14158) );
  NOR2X1 U12819 ( .A(n14162), .B(n14163), .Y(n14161) );
  OR2X1 U12820 ( .A(n14164), .B(n14165), .Y(n14163) );
  OAI21X1 U12821 ( .A(n12852), .B(n13958), .C(n14166), .Y(n14165) );
  AOI22X1 U12822 ( .A(n13960), .B(\regX[16][0] ), .C(n13961), .D(\regX[20][0] ), .Y(n14166) );
  AND2X1 U12823 ( .A(n14167), .B(n14168), .Y(n13961) );
  INVX1 U12824 ( .A(n14169), .Y(n13960) );
  NAND3X1 U12825 ( .A(n14168), .B(n14170), .C(n14171), .Y(n14169) );
  NAND2X1 U12826 ( .A(n14172), .B(n14167), .Y(n13958) );
  OAI21X1 U12827 ( .A(n12618), .B(n13962), .C(n14173), .Y(n14164) );
  AOI22X1 U12828 ( .A(n13964), .B(N1735), .C(n13965), .D(\regX[19][0] ), .Y(
        n14173) );
  AND2X1 U12829 ( .A(n14174), .B(n14175), .Y(n13965) );
  AND2X1 U12830 ( .A(n14172), .B(n14176), .Y(n13964) );
  NAND2X1 U12831 ( .A(n14177), .B(n14167), .Y(n13962) );
  INVX1 U12832 ( .A(\regX[13][0] ), .Y(n12618) );
  NAND3X1 U12833 ( .A(n14178), .B(n14179), .C(n14180), .Y(n14162) );
  AOI21X1 U12834 ( .A(n13969), .B(\regX[15][0] ), .C(n14181), .Y(n14180) );
  OAI22X1 U12835 ( .A(n12804), .B(n13971), .C(n12842), .D(n13972), .Y(n14181)
         );
  NAND2X1 U12836 ( .A(n14176), .B(n14174), .Y(n13972) );
  NAND2X1 U12837 ( .A(n14182), .B(n14183), .Y(n13971) );
  INVX1 U12838 ( .A(n14170), .Y(n14182) );
  AND2X1 U12839 ( .A(n14177), .B(n14176), .Y(n13969) );
  AOI22X1 U12840 ( .A(n13973), .B(\regX[18][0] ), .C(n13974), .D(\regX[21][0] ), .Y(n14179) );
  AND2X1 U12841 ( .A(n14167), .B(n14174), .Y(n13974) );
  AND2X1 U12842 ( .A(n14175), .B(n14168), .Y(n13973) );
  AOI22X1 U12843 ( .A(n13975), .B(\regX[22][0] ), .C(n13976), .D(\regX[17][0] ), .Y(n14178) );
  AND2X1 U12844 ( .A(n14171), .B(n14174), .Y(n13976) );
  NOR2X1 U12845 ( .A(n14184), .B(n14185), .Y(n14174) );
  AND2X1 U12846 ( .A(n14176), .B(n14168), .Y(n13975) );
  NOR2X1 U12847 ( .A(n14186), .B(n14184), .Y(n14168) );
  NOR2X1 U12848 ( .A(n14187), .B(n14188), .Y(n14160) );
  OAI21X1 U12849 ( .A(n12669), .B(n13979), .C(n14189), .Y(n14188) );
  AOI22X1 U12850 ( .A(n13981), .B(\regX[8][0] ), .C(n13982), .D(\regX[7][0] ), 
        .Y(n14189) );
  AND2X1 U12851 ( .A(n14190), .B(n14176), .Y(n13982) );
  INVX1 U12852 ( .A(n14191), .Y(n13981) );
  NAND3X1 U12853 ( .A(n14171), .B(n14184), .C(n14172), .Y(n14191) );
  NAND2X1 U12854 ( .A(n14192), .B(n14176), .Y(n13979) );
  NOR2X1 U12855 ( .A(n14193), .B(n14194), .Y(n14176) );
  OAI21X1 U12856 ( .A(n12771), .B(n13983), .C(n14195), .Y(n14187) );
  AOI22X1 U12857 ( .A(n13985), .B(\regX[11][0] ), .C(n13986), .D(N1615), .Y(
        n14195) );
  AND2X1 U12858 ( .A(n14172), .B(n14175), .Y(n13986) );
  NOR2X1 U12859 ( .A(n14170), .B(n14186), .Y(n14172) );
  AND2X1 U12860 ( .A(n14177), .B(n14175), .Y(n13985) );
  NAND2X1 U12861 ( .A(n14177), .B(n14171), .Y(n13983) );
  NOR2X1 U12862 ( .A(n14170), .B(n14185), .Y(n14177) );
  NOR2X1 U12863 ( .A(n14196), .B(n14197), .Y(n14159) );
  OAI21X1 U12864 ( .A(n12605), .B(n13989), .C(n14198), .Y(n14197) );
  AOI22X1 U12865 ( .A(n13991), .B(N1375), .C(n13992), .D(\regX[1][0] ), .Y(
        n14198) );
  AND2X1 U12866 ( .A(n14190), .B(n14171), .Y(n13992) );
  AND2X1 U12867 ( .A(n14192), .B(n14175), .Y(n13991) );
  NAND2X1 U12868 ( .A(n14192), .B(n14171), .Y(n13989) );
  NOR2X1 U12869 ( .A(n14199), .B(n14200), .Y(n14171) );
  INVX1 U12870 ( .A(\regX[0][0] ), .Y(n12605) );
  OAI21X1 U12871 ( .A(n12712), .B(n13993), .C(n14201), .Y(n14196) );
  AOI22X1 U12872 ( .A(n13995), .B(\regX[5][0] ), .C(n13996), .D(N1433), .Y(
        n14201) );
  AND2X1 U12873 ( .A(n14192), .B(n14167), .Y(n13996) );
  INVX1 U12874 ( .A(n14202), .Y(n14192) );
  NAND3X1 U12875 ( .A(n14170), .B(n14184), .C(n14185), .Y(n14202) );
  INVX1 U12876 ( .A(n14186), .Y(n14185) );
  AND2X1 U12877 ( .A(n14190), .B(n14167), .Y(n13995) );
  NOR2X1 U12878 ( .A(n14199), .B(n14193), .Y(n14167) );
  NAND2X1 U12879 ( .A(n14190), .B(n14175), .Y(n13993) );
  NOR2X1 U12880 ( .A(n14200), .B(n14194), .Y(n14175) );
  INVX1 U12881 ( .A(n14199), .Y(n14194) );
  INVX1 U12882 ( .A(n14203), .Y(n14190) );
  NAND3X1 U12883 ( .A(n14184), .B(n14186), .C(n14170), .Y(n14203) );
  INVX1 U12884 ( .A(n14183), .Y(n14184) );
  OAI21X1 U12885 ( .A(n12470), .B(n12869), .C(n14204), .Y(\U3/U91/Z_7 ) );
  OAI21X1 U12886 ( .A(n12470), .B(n12868), .C(n14204), .Y(\U3/U91/Z_6 ) );
  OAI21X1 U12887 ( .A(n12470), .B(n12867), .C(n14204), .Y(\U3/U91/Z_5 ) );
  OAI21X1 U12888 ( .A(n12470), .B(n12866), .C(n14204), .Y(\U3/U91/Z_4 ) );
  OAI21X1 U12889 ( .A(n12470), .B(n12865), .C(n14204), .Y(\U3/U91/Z_3 ) );
  OAI21X1 U12890 ( .A(n12470), .B(n12864), .C(n14204), .Y(\U3/U91/Z_2 ) );
  OAI21X1 U12891 ( .A(n12470), .B(n12863), .C(n14204), .Y(\U3/U91/Z_1 ) );
  NAND2X1 U12892 ( .A(dy[1]), .B(n15369), .Y(n14204) );
  OAI22X1 U12893 ( .A(n13921), .B(n12553), .C(n12470), .D(n12861), .Y(
        \U3/U91/Z_0 ) );
  NAND2X1 U12894 ( .A(n13921), .B(n12470), .Y(\U3/U90/Z_0 ) );
  OR2X1 U12895 ( .A(\U3/U122/Z_8 ), .B(n12476), .Y(\U3/U88/Z_9 ) );
  OAI21X1 U12896 ( .A(n12464), .B(n12970), .C(n12486), .Y(\U3/U88/Z_8 ) );
  OAI21X1 U12897 ( .A(n12470), .B(n12850), .C(n14205), .Y(\U3/U88/Z_7 ) );
  AOI21X1 U12898 ( .A(fGx[7]), .B(n12466), .C(n12476), .Y(n14205) );
  OAI21X1 U12899 ( .A(n12470), .B(n12849), .C(n14206), .Y(\U3/U88/Z_6 ) );
  AOI21X1 U12900 ( .A(fGx[6]), .B(n12466), .C(n12476), .Y(n14206) );
  OAI21X1 U12901 ( .A(n12470), .B(n12848), .C(n14207), .Y(\U3/U88/Z_5 ) );
  AOI21X1 U12902 ( .A(fGx[5]), .B(n12466), .C(n12476), .Y(n14207) );
  OAI21X1 U12903 ( .A(n12470), .B(n12847), .C(n14208), .Y(\U3/U88/Z_4 ) );
  AOI21X1 U12904 ( .A(fGx[4]), .B(n12466), .C(n12476), .Y(n14208) );
  OR2X1 U12905 ( .A(\U3/U122/Z_29 ), .B(n12476), .Y(\U3/U88/Z_30 ) );
  OAI21X1 U12906 ( .A(n12470), .B(n12846), .C(n14209), .Y(\U3/U88/Z_3 ) );
  AOI21X1 U12907 ( .A(fGx[3]), .B(n12466), .C(n12476), .Y(n14209) );
  OR2X1 U12908 ( .A(\U3/U122/Z_28 ), .B(n12476), .Y(\U3/U88/Z_29 ) );
  OR2X1 U12909 ( .A(\U3/U122/Z_27 ), .B(n12476), .Y(\U3/U88/Z_28 ) );
  OR2X1 U12910 ( .A(\U3/U122/Z_26 ), .B(n12476), .Y(\U3/U88/Z_27 ) );
  OR2X1 U12911 ( .A(\U3/U122/Z_25 ), .B(n12476), .Y(\U3/U88/Z_26 ) );
  OR2X1 U12912 ( .A(\U3/U122/Z_24 ), .B(n12476), .Y(\U3/U88/Z_25 ) );
  OR2X1 U12913 ( .A(\U3/U122/Z_23 ), .B(n12476), .Y(\U3/U88/Z_24 ) );
  OR2X1 U12914 ( .A(\U3/U122/Z_22 ), .B(n12476), .Y(\U3/U88/Z_23 ) );
  OR2X1 U12915 ( .A(\U3/U122/Z_21 ), .B(n12476), .Y(\U3/U88/Z_22 ) );
  OR2X1 U12916 ( .A(\U3/U122/Z_20 ), .B(n12476), .Y(\U3/U88/Z_21 ) );
  OR2X1 U12917 ( .A(\U3/U122/Z_19 ), .B(n12476), .Y(\U3/U88/Z_20 ) );
  OAI21X1 U12918 ( .A(n12470), .B(n12845), .C(n14210), .Y(\U3/U88/Z_2 ) );
  AOI21X1 U12919 ( .A(fGx[2]), .B(n12466), .C(n12476), .Y(n14210) );
  OR2X1 U12920 ( .A(\U3/U122/Z_18 ), .B(n12476), .Y(\U3/U88/Z_19 ) );
  OR2X1 U12921 ( .A(\U3/U122/Z_17 ), .B(n12476), .Y(\U3/U88/Z_18 ) );
  OR2X1 U12922 ( .A(\U3/U122/Z_16 ), .B(n12476), .Y(\U3/U88/Z_17 ) );
  OR2X1 U12923 ( .A(\U3/U122/Z_15 ), .B(n12476), .Y(\U3/U88/Z_16 ) );
  OR2X1 U12924 ( .A(\U3/U122/Z_14 ), .B(n12476), .Y(\U3/U88/Z_15 ) );
  OR2X1 U12925 ( .A(\U3/U122/Z_13 ), .B(n12476), .Y(\U3/U88/Z_14 ) );
  OR2X1 U12926 ( .A(\U3/U122/Z_12 ), .B(n12476), .Y(\U3/U88/Z_13 ) );
  OR2X1 U12927 ( .A(\U3/U122/Z_11 ), .B(n12476), .Y(\U3/U88/Z_12 ) );
  OR2X1 U12928 ( .A(\U3/U122/Z_10 ), .B(n12476), .Y(\U3/U88/Z_11 ) );
  OR2X1 U12929 ( .A(\U3/U122/Z_9 ), .B(n12476), .Y(\U3/U88/Z_10 ) );
  OAI21X1 U12930 ( .A(n12470), .B(n12844), .C(n14211), .Y(\U3/U88/Z_1 ) );
  AOI21X1 U12931 ( .A(fGx[1]), .B(n12466), .C(n12476), .Y(n14211) );
  OAI21X1 U12932 ( .A(n12470), .B(n12842), .C(n14212), .Y(\U3/U88/Z_0 ) );
  AOI21X1 U12933 ( .A(fGx[0]), .B(n12466), .C(n12476), .Y(n14212) );
  NOR2X1 U12934 ( .A(n12479), .B(n12860), .Y(\U3/U87/Z_7 ) );
  NOR2X1 U12935 ( .A(n12483), .B(n12859), .Y(\U3/U87/Z_6 ) );
  NOR2X1 U12936 ( .A(n12483), .B(n12858), .Y(\U3/U87/Z_5 ) );
  NOR2X1 U12937 ( .A(n12483), .B(n12857), .Y(\U3/U87/Z_4 ) );
  NOR2X1 U12938 ( .A(n12483), .B(n12856), .Y(\U3/U87/Z_3 ) );
  OAI21X1 U12939 ( .A(n12480), .B(n12855), .C(n12464), .Y(\U3/U87/Z_2 ) );
  OAI21X1 U12940 ( .A(n12481), .B(n12854), .C(n12470), .Y(\U3/U87/Z_1 ) );
  OAI21X1 U12941 ( .A(n12480), .B(n12852), .C(n14213), .Y(\U3/U87/Z_0 ) );
  NOR2X1 U12942 ( .A(n15370), .B(n12466), .Y(n14213) );
  OAI21X1 U12943 ( .A(n14214), .B(n13063), .C(n12488), .Y(\U3/U85/Z_9 ) );
  OAI21X1 U12944 ( .A(n14214), .B(n12970), .C(n12488), .Y(\U3/U85/Z_8 ) );
  OAI21X1 U12945 ( .A(n14214), .B(n14215), .C(n14216), .Y(\U3/U85/Z_7 ) );
  AOI21X1 U12946 ( .A(\regX[22][7] ), .B(n15370), .C(n12476), .Y(n14216) );
  OAI21X1 U12947 ( .A(n14214), .B(n14217), .C(n14218), .Y(\U3/U85/Z_6 ) );
  AOI21X1 U12948 ( .A(\regX[22][6] ), .B(n15370), .C(n12476), .Y(n14218) );
  OAI21X1 U12949 ( .A(n14214), .B(n14219), .C(n14220), .Y(\U3/U85/Z_5 ) );
  AOI21X1 U12950 ( .A(\regX[22][5] ), .B(n15370), .C(n12476), .Y(n14220) );
  OAI21X1 U12951 ( .A(n14214), .B(n14221), .C(n14222), .Y(\U3/U85/Z_4 ) );
  AOI21X1 U12952 ( .A(\regX[22][4] ), .B(n15370), .C(n12476), .Y(n14222) );
  OAI21X1 U12953 ( .A(n14214), .B(n13163), .C(n12488), .Y(\U3/U85/Z_31 ) );
  OAI21X1 U12954 ( .A(n14214), .B(n13159), .C(n12489), .Y(\U3/U85/Z_30 ) );
  OAI21X1 U12955 ( .A(n14214), .B(n14223), .C(n14224), .Y(\U3/U85/Z_3 ) );
  AOI21X1 U12956 ( .A(\regX[22][3] ), .B(n15370), .C(n12476), .Y(n14224) );
  OAI21X1 U12957 ( .A(n14214), .B(n13155), .C(n12488), .Y(\U3/U85/Z_29 ) );
  OAI21X1 U12958 ( .A(n14214), .B(n13151), .C(n12488), .Y(\U3/U85/Z_28 ) );
  OAI21X1 U12959 ( .A(n14214), .B(n13147), .C(n12488), .Y(\U3/U85/Z_27 ) );
  OAI21X1 U12960 ( .A(n14214), .B(n13143), .C(n12488), .Y(\U3/U85/Z_26 ) );
  OAI21X1 U12961 ( .A(n14214), .B(n13139), .C(n12488), .Y(\U3/U85/Z_25 ) );
  OAI21X1 U12962 ( .A(n14214), .B(n13135), .C(n12488), .Y(\U3/U85/Z_24 ) );
  OAI21X1 U12963 ( .A(n14214), .B(n13131), .C(n12488), .Y(\U3/U85/Z_23 ) );
  OAI21X1 U12964 ( .A(n14214), .B(n13127), .C(n12488), .Y(\U3/U85/Z_22 ) );
  OAI21X1 U12965 ( .A(n14214), .B(n13123), .C(n12487), .Y(\U3/U85/Z_21 ) );
  OAI21X1 U12966 ( .A(n14214), .B(n13119), .C(n12487), .Y(\U3/U85/Z_20 ) );
  OAI21X1 U12967 ( .A(n14214), .B(n14225), .C(n14226), .Y(\U3/U85/Z_2 ) );
  AOI21X1 U12968 ( .A(\regX[22][2] ), .B(n15370), .C(n12476), .Y(n14226) );
  OAI21X1 U12969 ( .A(n14214), .B(n13115), .C(n12487), .Y(\U3/U85/Z_19 ) );
  OAI21X1 U12970 ( .A(n14214), .B(n13111), .C(n12489), .Y(\U3/U85/Z_18 ) );
  OAI21X1 U12971 ( .A(n14214), .B(n13107), .C(n12487), .Y(\U3/U85/Z_17 ) );
  OAI21X1 U12972 ( .A(n14214), .B(n13103), .C(n12487), .Y(\U3/U85/Z_16 ) );
  OAI21X1 U12973 ( .A(n14214), .B(n13099), .C(n12487), .Y(\U3/U85/Z_15 ) );
  OAI21X1 U12974 ( .A(n14214), .B(n13095), .C(n12487), .Y(\U3/U85/Z_14 ) );
  OAI21X1 U12975 ( .A(n14214), .B(n13091), .C(n12487), .Y(\U3/U85/Z_13 ) );
  OAI21X1 U12976 ( .A(n14214), .B(n13087), .C(n12487), .Y(\U3/U85/Z_12 ) );
  OAI21X1 U12977 ( .A(n14214), .B(n13083), .C(n12486), .Y(\U3/U85/Z_11 ) );
  OAI21X1 U12978 ( .A(n14214), .B(n13079), .C(n12487), .Y(\U3/U85/Z_10 ) );
  OAI21X1 U12979 ( .A(n14214), .B(n14227), .C(n14228), .Y(\U3/U85/Z_1 ) );
  AOI21X1 U12980 ( .A(\regX[22][1] ), .B(n15370), .C(n12476), .Y(n14228) );
  OAI22X1 U12981 ( .A(n14214), .B(n14229), .C(n12470), .D(n12832), .Y(
        \U3/U85/Z_0 ) );
  OAI21X1 U12982 ( .A(n12480), .B(n12899), .C(n14214), .Y(\U3/U84/Z_7 ) );
  OAI21X1 U12983 ( .A(n12480), .B(n12898), .C(n14214), .Y(\U3/U84/Z_6 ) );
  OAI21X1 U12984 ( .A(n12481), .B(n12897), .C(n14214), .Y(\U3/U84/Z_5 ) );
  OAI21X1 U12985 ( .A(n12480), .B(n12896), .C(n14214), .Y(\U3/U84/Z_4 ) );
  OAI21X1 U12986 ( .A(n12481), .B(n12895), .C(n14214), .Y(\U3/U84/Z_3 ) );
  INVX1 U12987 ( .A(\regX[11][3] ), .Y(n12895) );
  OAI21X1 U12988 ( .A(n12481), .B(n12894), .C(n12470), .Y(\U3/U84/Z_2 ) );
  INVX1 U12989 ( .A(\regX[11][2] ), .Y(n12894) );
  OAI21X1 U12990 ( .A(n12481), .B(n12893), .C(n14214), .Y(\U3/U84/Z_1 ) );
  INVX1 U12991 ( .A(\regX[11][1] ), .Y(n12893) );
  OAI21X1 U12992 ( .A(n12482), .B(n12891), .C(n14214), .Y(\U3/U84/Z_0 ) );
  INVX1 U12993 ( .A(\regX[11][0] ), .Y(n12891) );
  OAI21X1 U12994 ( .A(n13892), .B(n13063), .C(n14230), .Y(\U3/U82/Z_9 ) );
  AOI22X1 U12995 ( .A(n12475), .B(Gy[9]), .C(N2245), .D(n12471), .Y(n14230) );
  OAI21X1 U12996 ( .A(n13892), .B(n12970), .C(n14231), .Y(\U3/U82/Z_8 ) );
  AOI22X1 U12997 ( .A(n12475), .B(Gy[8]), .C(N2244), .D(n12471), .Y(n14231) );
  OAI21X1 U12998 ( .A(n13892), .B(n14215), .C(n14232), .Y(\U3/U82/Z_7 ) );
  AOI22X1 U12999 ( .A(n12475), .B(Gy[7]), .C(N2243), .D(n12471), .Y(n14232) );
  OAI21X1 U13000 ( .A(n13892), .B(n14217), .C(n14233), .Y(\U3/U82/Z_6 ) );
  AOI22X1 U13001 ( .A(n12475), .B(Gy[6]), .C(N2242), .D(n12471), .Y(n14233) );
  OAI21X1 U13002 ( .A(n13892), .B(n14219), .C(n14234), .Y(\U3/U82/Z_5 ) );
  AOI22X1 U13003 ( .A(n12475), .B(Gy[5]), .C(N2241), .D(n12471), .Y(n14234) );
  OAI21X1 U13004 ( .A(n13892), .B(n14221), .C(n14235), .Y(\U3/U82/Z_4 ) );
  AOI22X1 U13005 ( .A(n12475), .B(Gy[4]), .C(N2240), .D(n12471), .Y(n14235) );
  OAI21X1 U13006 ( .A(n13892), .B(n13163), .C(n14236), .Y(\U3/U82/Z_31 ) );
  AOI21X1 U13007 ( .A(N2267), .B(n12471), .C(n12475), .Y(n14236) );
  OAI21X1 U13008 ( .A(n13892), .B(n13159), .C(n14237), .Y(\U3/U82/Z_30 ) );
  AOI22X1 U13009 ( .A(n12475), .B(Gy[30]), .C(N2266), .D(n12471), .Y(n14237)
         );
  OAI21X1 U13010 ( .A(n13892), .B(n14223), .C(n14238), .Y(\U3/U82/Z_3 ) );
  AOI22X1 U13011 ( .A(n12475), .B(Gy[3]), .C(N2239), .D(n12471), .Y(n14238) );
  OAI21X1 U13012 ( .A(n13892), .B(n13155), .C(n14239), .Y(\U3/U82/Z_29 ) );
  AOI22X1 U13013 ( .A(n12475), .B(Gy[29]), .C(N2265), .D(n12471), .Y(n14239)
         );
  OAI21X1 U13014 ( .A(n13892), .B(n13151), .C(n14240), .Y(\U3/U82/Z_28 ) );
  AOI22X1 U13015 ( .A(n12475), .B(Gy[28]), .C(N2264), .D(n12471), .Y(n14240)
         );
  OAI21X1 U13016 ( .A(n13892), .B(n13147), .C(n14241), .Y(\U3/U82/Z_27 ) );
  AOI22X1 U13017 ( .A(n12475), .B(Gy[27]), .C(N2263), .D(n12471), .Y(n14241)
         );
  OAI21X1 U13018 ( .A(n13892), .B(n13143), .C(n14242), .Y(\U3/U82/Z_26 ) );
  AOI22X1 U13019 ( .A(n12475), .B(Gy[26]), .C(N2262), .D(n12471), .Y(n14242)
         );
  OAI21X1 U13020 ( .A(n13892), .B(n13139), .C(n14243), .Y(\U3/U82/Z_25 ) );
  AOI22X1 U13021 ( .A(n12475), .B(Gy[25]), .C(N2261), .D(n12471), .Y(n14243)
         );
  OAI21X1 U13022 ( .A(n13892), .B(n13135), .C(n14244), .Y(\U3/U82/Z_24 ) );
  AOI22X1 U13023 ( .A(n12475), .B(Gy[24]), .C(N2260), .D(n12471), .Y(n14244)
         );
  OAI21X1 U13024 ( .A(n13892), .B(n13131), .C(n14245), .Y(\U3/U82/Z_23 ) );
  AOI22X1 U13025 ( .A(n12475), .B(Gy[23]), .C(N2259), .D(n12471), .Y(n14245)
         );
  OAI21X1 U13026 ( .A(n13892), .B(n13127), .C(n14246), .Y(\U3/U82/Z_22 ) );
  AOI22X1 U13027 ( .A(n12475), .B(Gy[22]), .C(N2258), .D(n12471), .Y(n14246)
         );
  OAI21X1 U13028 ( .A(n13892), .B(n13123), .C(n14247), .Y(\U3/U82/Z_21 ) );
  AOI22X1 U13029 ( .A(n12475), .B(Gy[21]), .C(N2257), .D(n12471), .Y(n14247)
         );
  OAI21X1 U13030 ( .A(n13892), .B(n13119), .C(n14248), .Y(\U3/U82/Z_20 ) );
  AOI22X1 U13031 ( .A(n12475), .B(Gy[20]), .C(N2256), .D(n12471), .Y(n14248)
         );
  OAI21X1 U13032 ( .A(n13892), .B(n14225), .C(n14249), .Y(\U3/U82/Z_2 ) );
  AOI22X1 U13033 ( .A(n12475), .B(Gy[2]), .C(N2238), .D(n12471), .Y(n14249) );
  OAI21X1 U13034 ( .A(n13892), .B(n13115), .C(n14250), .Y(\U3/U82/Z_19 ) );
  AOI22X1 U13035 ( .A(n12475), .B(Gy[19]), .C(N2255), .D(n12471), .Y(n14250)
         );
  OAI21X1 U13036 ( .A(n13892), .B(n13111), .C(n14251), .Y(\U3/U82/Z_18 ) );
  AOI22X1 U13037 ( .A(n12475), .B(Gy[18]), .C(N2254), .D(n12471), .Y(n14251)
         );
  OAI21X1 U13038 ( .A(n13892), .B(n13107), .C(n14252), .Y(\U3/U82/Z_17 ) );
  AOI22X1 U13039 ( .A(n12475), .B(Gy[17]), .C(N2253), .D(n12471), .Y(n14252)
         );
  OAI21X1 U13040 ( .A(n13892), .B(n13103), .C(n14253), .Y(\U3/U82/Z_16 ) );
  AOI22X1 U13041 ( .A(n12475), .B(Gy[16]), .C(N2252), .D(n12471), .Y(n14253)
         );
  OAI21X1 U13042 ( .A(n13892), .B(n13099), .C(n14254), .Y(\U3/U82/Z_15 ) );
  AOI22X1 U13043 ( .A(n12475), .B(Gy[15]), .C(N2251), .D(n12471), .Y(n14254)
         );
  OAI21X1 U13044 ( .A(n13892), .B(n13095), .C(n14255), .Y(\U3/U82/Z_14 ) );
  AOI22X1 U13045 ( .A(n12475), .B(Gy[14]), .C(N2250), .D(n12471), .Y(n14255)
         );
  OAI21X1 U13046 ( .A(n13892), .B(n13091), .C(n14256), .Y(\U3/U82/Z_13 ) );
  AOI22X1 U13047 ( .A(n12475), .B(Gy[13]), .C(N2249), .D(n12471), .Y(n14256)
         );
  OAI21X1 U13048 ( .A(n13892), .B(n13087), .C(n14257), .Y(\U3/U82/Z_12 ) );
  AOI22X1 U13049 ( .A(n12475), .B(Gy[12]), .C(N2248), .D(n12471), .Y(n14257)
         );
  OAI21X1 U13050 ( .A(n13892), .B(n13083), .C(n14258), .Y(\U3/U82/Z_11 ) );
  AOI22X1 U13051 ( .A(n12475), .B(Gy[11]), .C(N2247), .D(n12471), .Y(n14258)
         );
  OAI21X1 U13052 ( .A(n13892), .B(n13079), .C(n14259), .Y(\U3/U82/Z_10 ) );
  AOI22X1 U13053 ( .A(n12475), .B(Gy[10]), .C(N2246), .D(n12471), .Y(n14259)
         );
  OAI21X1 U13054 ( .A(n13892), .B(n14227), .C(n14260), .Y(\U3/U82/Z_1 ) );
  AOI22X1 U13055 ( .A(n12475), .B(Gy[1]), .C(N2237), .D(n12471), .Y(n14260) );
  OAI21X1 U13056 ( .A(n13892), .B(n14229), .C(n14261), .Y(\U3/U82/Z_0 ) );
  AOI22X1 U13057 ( .A(n12475), .B(Gy[0]), .C(N2236), .D(n12471), .Y(n14261) );
  INVX1 U13058 ( .A(fGx[0]), .Y(n14229) );
  NOR2X1 U13059 ( .A(n12462), .B(n12860), .Y(\U3/U81/Z_7 ) );
  NOR2X1 U13060 ( .A(n12462), .B(n12859), .Y(\U3/U81/Z_6 ) );
  NOR2X1 U13061 ( .A(n12462), .B(n12858), .Y(\U3/U81/Z_5 ) );
  NOR2X1 U13062 ( .A(n12462), .B(n12857), .Y(\U3/U81/Z_4 ) );
  NOR2X1 U13063 ( .A(n12462), .B(n12856), .Y(\U3/U81/Z_3 ) );
  NOR2X1 U13064 ( .A(n12462), .B(n12855), .Y(\U3/U81/Z_2 ) );
  NOR2X1 U13065 ( .A(n12462), .B(n12854), .Y(\U3/U81/Z_1 ) );
  NOR2X1 U13066 ( .A(n12462), .B(n12852), .Y(\U3/U81/Z_0 ) );
  OAI21X1 U13067 ( .A(n13893), .B(n13061), .C(n14262), .Y(\U3/U79/Z_9 ) );
  NAND2X1 U13068 ( .A(N2277), .B(n12471), .Y(n14262) );
  INVX1 U13069 ( .A(Gx[9]), .Y(n13061) );
  OAI21X1 U13070 ( .A(n13893), .B(n13059), .C(n14263), .Y(\U3/U79/Z_8 ) );
  NAND2X1 U13071 ( .A(N2276), .B(n12471), .Y(n14263) );
  INVX1 U13072 ( .A(Gx[8]), .Y(n13059) );
  OAI21X1 U13073 ( .A(n13893), .B(n13055), .C(n14264), .Y(\U3/U79/Z_7 ) );
  NAND2X1 U13074 ( .A(N2275), .B(n12471), .Y(n14264) );
  INVX1 U13075 ( .A(Gx[7]), .Y(n13055) );
  OAI21X1 U13076 ( .A(n13893), .B(n13052), .C(n14265), .Y(\U3/U79/Z_6 ) );
  NAND2X1 U13077 ( .A(N2274), .B(n12471), .Y(n14265) );
  INVX1 U13078 ( .A(Gx[6]), .Y(n13052) );
  OAI21X1 U13079 ( .A(n13893), .B(n13049), .C(n14266), .Y(\U3/U79/Z_5 ) );
  NAND2X1 U13080 ( .A(N2273), .B(n12471), .Y(n14266) );
  INVX1 U13081 ( .A(Gx[5]), .Y(n13049) );
  OAI21X1 U13082 ( .A(n13893), .B(n13046), .C(n14267), .Y(\U3/U79/Z_4 ) );
  NAND2X1 U13083 ( .A(N2272), .B(n12471), .Y(n14267) );
  INVX1 U13084 ( .A(Gx[4]), .Y(n13046) );
  OAI21X1 U13085 ( .A(n13893), .B(n13161), .C(n14268), .Y(\U3/U79/Z_31 ) );
  NAND2X1 U13086 ( .A(N2299), .B(n12471), .Y(n14268) );
  INVX1 U13087 ( .A(Gx[31]), .Y(n13161) );
  OAI21X1 U13088 ( .A(n13893), .B(n13157), .C(n14269), .Y(\U3/U79/Z_30 ) );
  NAND2X1 U13089 ( .A(N2298), .B(n12471), .Y(n14269) );
  INVX1 U13090 ( .A(Gx[30]), .Y(n13157) );
  OAI21X1 U13091 ( .A(n13893), .B(n13043), .C(n14270), .Y(\U3/U79/Z_3 ) );
  NAND2X1 U13092 ( .A(N2271), .B(n12471), .Y(n14270) );
  INVX1 U13093 ( .A(Gx[3]), .Y(n13043) );
  OAI21X1 U13094 ( .A(n13893), .B(n13153), .C(n14271), .Y(\U3/U79/Z_29 ) );
  NAND2X1 U13095 ( .A(N2297), .B(n12471), .Y(n14271) );
  INVX1 U13096 ( .A(Gx[29]), .Y(n13153) );
  OAI21X1 U13097 ( .A(n13893), .B(n13149), .C(n14272), .Y(\U3/U79/Z_28 ) );
  NAND2X1 U13098 ( .A(N2296), .B(n12471), .Y(n14272) );
  INVX1 U13099 ( .A(Gx[28]), .Y(n13149) );
  OAI21X1 U13100 ( .A(n13893), .B(n13145), .C(n14273), .Y(\U3/U79/Z_27 ) );
  NAND2X1 U13101 ( .A(N2295), .B(n12471), .Y(n14273) );
  INVX1 U13102 ( .A(Gx[27]), .Y(n13145) );
  OAI21X1 U13103 ( .A(n13893), .B(n13141), .C(n14274), .Y(\U3/U79/Z_26 ) );
  NAND2X1 U13104 ( .A(N2294), .B(n12471), .Y(n14274) );
  INVX1 U13105 ( .A(Gx[26]), .Y(n13141) );
  OAI21X1 U13106 ( .A(n13893), .B(n13137), .C(n14275), .Y(\U3/U79/Z_25 ) );
  NAND2X1 U13107 ( .A(N2293), .B(n12471), .Y(n14275) );
  INVX1 U13108 ( .A(Gx[25]), .Y(n13137) );
  OAI21X1 U13109 ( .A(n13893), .B(n13133), .C(n14276), .Y(\U3/U79/Z_24 ) );
  NAND2X1 U13110 ( .A(N2292), .B(n12471), .Y(n14276) );
  INVX1 U13111 ( .A(Gx[24]), .Y(n13133) );
  OAI21X1 U13112 ( .A(n13893), .B(n13129), .C(n14277), .Y(\U3/U79/Z_23 ) );
  NAND2X1 U13113 ( .A(N2291), .B(n12471), .Y(n14277) );
  INVX1 U13114 ( .A(Gx[23]), .Y(n13129) );
  OAI21X1 U13115 ( .A(n13893), .B(n13125), .C(n14278), .Y(\U3/U79/Z_22 ) );
  NAND2X1 U13116 ( .A(N2290), .B(n12471), .Y(n14278) );
  INVX1 U13117 ( .A(Gx[22]), .Y(n13125) );
  OAI21X1 U13118 ( .A(n13893), .B(n13121), .C(n14279), .Y(\U3/U79/Z_21 ) );
  NAND2X1 U13119 ( .A(N2289), .B(n12471), .Y(n14279) );
  INVX1 U13120 ( .A(Gx[21]), .Y(n13121) );
  OAI21X1 U13121 ( .A(n13893), .B(n13117), .C(n14280), .Y(\U3/U79/Z_20 ) );
  NAND2X1 U13122 ( .A(N2288), .B(n12471), .Y(n14280) );
  INVX1 U13123 ( .A(Gx[20]), .Y(n13117) );
  OAI21X1 U13124 ( .A(n13893), .B(n13040), .C(n14281), .Y(\U3/U79/Z_2 ) );
  NAND2X1 U13125 ( .A(N2270), .B(n12471), .Y(n14281) );
  INVX1 U13126 ( .A(Gx[2]), .Y(n13040) );
  OAI21X1 U13127 ( .A(n13893), .B(n13113), .C(n14282), .Y(\U3/U79/Z_19 ) );
  NAND2X1 U13128 ( .A(N2287), .B(n12471), .Y(n14282) );
  INVX1 U13129 ( .A(Gx[19]), .Y(n13113) );
  OAI21X1 U13130 ( .A(n13893), .B(n13109), .C(n14283), .Y(\U3/U79/Z_18 ) );
  NAND2X1 U13131 ( .A(N2286), .B(n12471), .Y(n14283) );
  INVX1 U13132 ( .A(Gx[18]), .Y(n13109) );
  OAI21X1 U13133 ( .A(n13893), .B(n13105), .C(n14284), .Y(\U3/U79/Z_17 ) );
  NAND2X1 U13134 ( .A(N2285), .B(n12471), .Y(n14284) );
  INVX1 U13135 ( .A(Gx[17]), .Y(n13105) );
  OAI21X1 U13136 ( .A(n13893), .B(n13101), .C(n14285), .Y(\U3/U79/Z_16 ) );
  NAND2X1 U13137 ( .A(N2284), .B(n12471), .Y(n14285) );
  INVX1 U13138 ( .A(Gx[16]), .Y(n13101) );
  OAI21X1 U13139 ( .A(n13893), .B(n13097), .C(n14286), .Y(\U3/U79/Z_15 ) );
  NAND2X1 U13140 ( .A(N2283), .B(n12471), .Y(n14286) );
  INVX1 U13141 ( .A(Gx[15]), .Y(n13097) );
  OAI21X1 U13142 ( .A(n13893), .B(n13093), .C(n14287), .Y(\U3/U79/Z_14 ) );
  NAND2X1 U13143 ( .A(N2282), .B(n12471), .Y(n14287) );
  INVX1 U13144 ( .A(Gx[14]), .Y(n13093) );
  OAI21X1 U13145 ( .A(n13893), .B(n13089), .C(n14288), .Y(\U3/U79/Z_13 ) );
  NAND2X1 U13146 ( .A(N2281), .B(n12471), .Y(n14288) );
  INVX1 U13147 ( .A(Gx[13]), .Y(n13089) );
  OAI21X1 U13148 ( .A(n13893), .B(n13085), .C(n14289), .Y(\U3/U79/Z_12 ) );
  NAND2X1 U13149 ( .A(N2280), .B(n12471), .Y(n14289) );
  INVX1 U13150 ( .A(Gx[12]), .Y(n13085) );
  OAI21X1 U13151 ( .A(n13893), .B(n13081), .C(n14290), .Y(\U3/U79/Z_11 ) );
  NAND2X1 U13152 ( .A(N2279), .B(n12471), .Y(n14290) );
  INVX1 U13153 ( .A(Gx[11]), .Y(n13081) );
  OAI21X1 U13154 ( .A(n13893), .B(n13065), .C(n14291), .Y(\U3/U79/Z_10 ) );
  NAND2X1 U13155 ( .A(N2278), .B(n12471), .Y(n14291) );
  INVX1 U13156 ( .A(Gx[10]), .Y(n13065) );
  OAI21X1 U13157 ( .A(n13893), .B(n13037), .C(n14292), .Y(\U3/U79/Z_1 ) );
  NAND2X1 U13158 ( .A(N2269), .B(n12471), .Y(n14292) );
  INVX1 U13159 ( .A(Gx[1]), .Y(n13037) );
  OAI21X1 U13160 ( .A(n13893), .B(n13033), .C(n14293), .Y(\U3/U79/Z_0 ) );
  NAND2X1 U13161 ( .A(N2268), .B(n12471), .Y(n14293) );
  INVX1 U13162 ( .A(Gx[0]), .Y(n13033) );
  NOR2X1 U13163 ( .A(n13165), .B(IntSignal[0]), .Y(n15363) );
  NOR2X1 U13164 ( .A(n12462), .B(n14294), .Y(\U3/U78/Z_9 ) );
  AND2X1 U13165 ( .A(n12471), .B(N2753), .Y(\U3/U78/Z_8 ) );
  AND2X1 U13166 ( .A(n12471), .B(N2752), .Y(\U3/U78/Z_7 ) );
  AND2X1 U13167 ( .A(n12471), .B(N2751), .Y(\U3/U78/Z_6 ) );
  AND2X1 U13168 ( .A(n12471), .B(N2750), .Y(\U3/U78/Z_5 ) );
  NOR2X1 U13169 ( .A(n12462), .B(n14295), .Y(\U3/U78/Z_4 ) );
  NOR2X1 U13170 ( .A(n12462), .B(n13032), .Y(\U3/U78/Z_31 ) );
  NOR2X1 U13171 ( .A(n12462), .B(n14296), .Y(\U3/U78/Z_30 ) );
  NOR2X1 U13172 ( .A(n12462), .B(n14297), .Y(\U3/U78/Z_3 ) );
  NOR2X1 U13173 ( .A(n12462), .B(n14298), .Y(\U3/U78/Z_29 ) );
  NOR2X1 U13174 ( .A(n12462), .B(n14299), .Y(\U3/U78/Z_28 ) );
  NOR2X1 U13175 ( .A(n12462), .B(n14300), .Y(\U3/U78/Z_27 ) );
  NOR2X1 U13176 ( .A(n12462), .B(n14301), .Y(\U3/U78/Z_26 ) );
  NOR2X1 U13177 ( .A(n12462), .B(n14302), .Y(\U3/U78/Z_25 ) );
  NOR2X1 U13178 ( .A(n12462), .B(n14303), .Y(\U3/U78/Z_24 ) );
  NOR2X1 U13179 ( .A(n12462), .B(n14304), .Y(\U3/U78/Z_23 ) );
  NOR2X1 U13180 ( .A(n12462), .B(n14305), .Y(\U3/U78/Z_22 ) );
  NOR2X1 U13181 ( .A(n12462), .B(n14306), .Y(\U3/U78/Z_21 ) );
  NOR2X1 U13182 ( .A(n12462), .B(n14307), .Y(\U3/U78/Z_20 ) );
  NOR2X1 U13183 ( .A(n12462), .B(n14308), .Y(\U3/U78/Z_2 ) );
  NOR2X1 U13184 ( .A(n12462), .B(n14309), .Y(\U3/U78/Z_19 ) );
  NOR2X1 U13185 ( .A(n12462), .B(n14310), .Y(\U3/U78/Z_18 ) );
  NOR2X1 U13186 ( .A(n12462), .B(n14311), .Y(\U3/U78/Z_17 ) );
  NOR2X1 U13187 ( .A(n12462), .B(n14312), .Y(\U3/U78/Z_16 ) );
  NOR2X1 U13188 ( .A(n12462), .B(n14313), .Y(\U3/U78/Z_15 ) );
  NOR2X1 U13189 ( .A(n12462), .B(n14314), .Y(\U3/U78/Z_14 ) );
  NOR2X1 U13190 ( .A(n12462), .B(n14315), .Y(\U3/U78/Z_13 ) );
  NOR2X1 U13191 ( .A(n12462), .B(n14316), .Y(\U3/U78/Z_12 ) );
  NOR2X1 U13192 ( .A(n12462), .B(n14317), .Y(\U3/U78/Z_11 ) );
  NOR2X1 U13193 ( .A(n12462), .B(n14318), .Y(\U3/U78/Z_10 ) );
  NOR2X1 U13194 ( .A(n12462), .B(n14319), .Y(\U3/U78/Z_1 ) );
  AND2X1 U13195 ( .A(n12471), .B(N2648), .Y(\U3/U78/Z_0 ) );
  AND2X1 U13196 ( .A(\U3/U77/DATA2_31 ), .B(n12477), .Y(\U3/U77/Z_31 ) );
  AND2X1 U13197 ( .A(\U3/U77/DATA2_30 ), .B(n12477), .Y(\U3/U77/Z_30 ) );
  AND2X1 U13198 ( .A(\U3/U77/DATA2_29 ), .B(n12477), .Y(\U3/U77/Z_29 ) );
  AND2X1 U13199 ( .A(\U3/U77/DATA2_28 ), .B(n12477), .Y(\U3/U77/Z_28 ) );
  AND2X1 U13200 ( .A(\U3/U77/DATA2_27 ), .B(n12477), .Y(\U3/U77/Z_27 ) );
  AND2X1 U13201 ( .A(\U3/U77/DATA2_26 ), .B(n12477), .Y(\U3/U77/Z_26 ) );
  AND2X1 U13202 ( .A(\U3/U77/DATA2_25 ), .B(n12477), .Y(\U3/U77/Z_25 ) );
  AND2X1 U13203 ( .A(\U3/U77/DATA2_24 ), .B(n12477), .Y(\U3/U77/Z_24 ) );
  AND2X1 U13204 ( .A(\U3/U77/DATA2_23 ), .B(n12477), .Y(\U3/U77/Z_23 ) );
  AND2X1 U13205 ( .A(\U3/U77/DATA2_22 ), .B(n12477), .Y(\U3/U77/Z_22 ) );
  AND2X1 U13206 ( .A(\U3/U77/DATA2_21 ), .B(n12477), .Y(\U3/U77/Z_21 ) );
  AND2X1 U13207 ( .A(\U3/U77/DATA2_20 ), .B(n12477), .Y(\U3/U77/Z_20 ) );
  AND2X1 U13208 ( .A(\U3/U77/DATA2_19 ), .B(n12477), .Y(\U3/U77/Z_19 ) );
  AND2X1 U13209 ( .A(\U3/U77/DATA2_18 ), .B(n12477), .Y(\U3/U77/Z_18 ) );
  AND2X1 U13210 ( .A(\U3/U77/DATA2_17 ), .B(n12477), .Y(\U3/U77/Z_17 ) );
  AND2X1 U13211 ( .A(\U3/U77/DATA2_16 ), .B(n12477), .Y(\U3/U77/Z_16 ) );
  AND2X1 U13212 ( .A(\U3/U77/DATA2_15 ), .B(n12477), .Y(\U3/U77/Z_15 ) );
  AND2X1 U13213 ( .A(N2399), .B(n15370), .Y(\U3/U76/Z_14 ) );
  AND2X1 U13214 ( .A(N2398), .B(n15370), .Y(\U3/U76/Z_13 ) );
  AND2X1 U13215 ( .A(N2397), .B(n15370), .Y(\U3/U76/Z_12 ) );
  AND2X1 U13216 ( .A(N2396), .B(n15370), .Y(\U3/U76/Z_11 ) );
  AND2X1 U13217 ( .A(N2395), .B(n15370), .Y(\U3/U76/Z_10 ) );
  AND2X1 U13218 ( .A(N2117), .B(n15370), .Y(\U3/U75/Z_9 ) );
  AND2X1 U13219 ( .A(N2116), .B(n15370), .Y(\U3/U75/Z_8 ) );
  OAI21X1 U13220 ( .A(n12482), .B(n12709), .C(n14320), .Y(\U3/U75/Z_7 ) );
  NAND2X1 U13221 ( .A(N2115), .B(n15370), .Y(n14320) );
  OAI21X1 U13222 ( .A(n12482), .B(n12708), .C(n14321), .Y(\U3/U75/Z_6 ) );
  NAND2X1 U13223 ( .A(N2114), .B(n15370), .Y(n14321) );
  OAI21X1 U13224 ( .A(n12483), .B(n12707), .C(n14322), .Y(\U3/U75/Z_5 ) );
  NAND2X1 U13225 ( .A(N2113), .B(n15370), .Y(n14322) );
  OAI21X1 U13226 ( .A(n12482), .B(n12706), .C(n14323), .Y(\U3/U75/Z_4 ) );
  NAND2X1 U13227 ( .A(N2112), .B(n15370), .Y(n14323) );
  OAI21X1 U13228 ( .A(n12483), .B(n12705), .C(n14324), .Y(\U3/U75/Z_3 ) );
  NAND2X1 U13229 ( .A(N2111), .B(n15370), .Y(n14324) );
  OAI21X1 U13230 ( .A(n12483), .B(n12704), .C(n14325), .Y(\U3/U75/Z_2 ) );
  NAND2X1 U13231 ( .A(N2110), .B(n15370), .Y(n14325) );
  AND2X1 U13232 ( .A(N2122), .B(n15370), .Y(\U3/U75/Z_14 ) );
  AND2X1 U13233 ( .A(N2121), .B(n15370), .Y(\U3/U75/Z_13 ) );
  AND2X1 U13234 ( .A(N2120), .B(n15370), .Y(\U3/U75/Z_12 ) );
  AND2X1 U13235 ( .A(N2119), .B(n15370), .Y(\U3/U75/Z_11 ) );
  AND2X1 U13236 ( .A(N2118), .B(n15370), .Y(\U3/U75/Z_10 ) );
  OAI21X1 U13237 ( .A(n12483), .B(n12703), .C(n14326), .Y(\U3/U75/Z_1 ) );
  NAND2X1 U13238 ( .A(N2109), .B(n15370), .Y(n14326) );
  OAI21X1 U13239 ( .A(n12483), .B(n12701), .C(n14327), .Y(\U3/U75/Z_0 ) );
  NAND2X1 U13240 ( .A(N2108), .B(n15370), .Y(n14327) );
  AND2X1 U13241 ( .A(n12477), .B(N2267), .Y(\U3/U74/Z_31 ) );
  AND2X1 U13242 ( .A(n12477), .B(N2266), .Y(\U3/U74/Z_30 ) );
  AND2X1 U13243 ( .A(n12477), .B(N2265), .Y(\U3/U74/Z_29 ) );
  AND2X1 U13244 ( .A(n12476), .B(N2264), .Y(\U3/U74/Z_28 ) );
  AND2X1 U13245 ( .A(n12476), .B(N2263), .Y(\U3/U74/Z_27 ) );
  AND2X1 U13246 ( .A(n12476), .B(N2262), .Y(\U3/U74/Z_26 ) );
  AND2X1 U13247 ( .A(n12476), .B(N2261), .Y(\U3/U74/Z_25 ) );
  AND2X1 U13248 ( .A(n12476), .B(N2260), .Y(\U3/U74/Z_24 ) );
  AND2X1 U13249 ( .A(n12476), .B(N2259), .Y(\U3/U74/Z_23 ) );
  AND2X1 U13250 ( .A(n12476), .B(N2258), .Y(\U3/U74/Z_22 ) );
  AND2X1 U13251 ( .A(n12476), .B(N2257), .Y(\U3/U74/Z_21 ) );
  AND2X1 U13252 ( .A(n12476), .B(N2256), .Y(\U3/U74/Z_20 ) );
  AND2X1 U13253 ( .A(n12476), .B(N2255), .Y(\U3/U74/Z_19 ) );
  AND2X1 U13254 ( .A(n12476), .B(N2254), .Y(\U3/U74/Z_18 ) );
  AND2X1 U13255 ( .A(n12476), .B(N2253), .Y(\U3/U74/Z_17 ) );
  AND2X1 U13256 ( .A(n12476), .B(N2252), .Y(\U3/U74/Z_16 ) );
  AND2X1 U13257 ( .A(n12476), .B(N2251), .Y(\U3/U74/Z_15 ) );
  NOR2X1 U13258 ( .A(n12484), .B(n13926), .Y(\U3/U73/Z_31 ) );
  INVX1 U13259 ( .A(N2911), .Y(n13926) );
  NOR2X1 U13260 ( .A(n12484), .B(n13928), .Y(\U3/U73/Z_30 ) );
  INVX1 U13261 ( .A(N2910), .Y(n13928) );
  NOR2X1 U13262 ( .A(n12484), .B(n13929), .Y(\U3/U73/Z_29 ) );
  INVX1 U13263 ( .A(N2909), .Y(n13929) );
  NOR2X1 U13264 ( .A(n12484), .B(n13930), .Y(\U3/U73/Z_28 ) );
  INVX1 U13265 ( .A(N2908), .Y(n13930) );
  NOR2X1 U13266 ( .A(n12484), .B(n13931), .Y(\U3/U73/Z_27 ) );
  INVX1 U13267 ( .A(N2907), .Y(n13931) );
  NOR2X1 U13268 ( .A(n12484), .B(n13932), .Y(\U3/U73/Z_26 ) );
  INVX1 U13269 ( .A(N2906), .Y(n13932) );
  NOR2X1 U13270 ( .A(n12484), .B(n13933), .Y(\U3/U73/Z_25 ) );
  INVX1 U13271 ( .A(N2905), .Y(n13933) );
  NOR2X1 U13272 ( .A(n12484), .B(n13934), .Y(\U3/U73/Z_24 ) );
  INVX1 U13273 ( .A(N2904), .Y(n13934) );
  NOR2X1 U13274 ( .A(n12484), .B(n13935), .Y(\U3/U73/Z_23 ) );
  INVX1 U13275 ( .A(N2903), .Y(n13935) );
  NOR2X1 U13276 ( .A(n12485), .B(n13936), .Y(\U3/U73/Z_22 ) );
  INVX1 U13277 ( .A(N2902), .Y(n13936) );
  NOR2X1 U13278 ( .A(n12485), .B(n13937), .Y(\U3/U73/Z_21 ) );
  INVX1 U13279 ( .A(N2901), .Y(n13937) );
  NOR2X1 U13280 ( .A(n12485), .B(n13939), .Y(\U3/U73/Z_20 ) );
  INVX1 U13281 ( .A(N2900), .Y(n13939) );
  NOR2X1 U13282 ( .A(n12485), .B(n13940), .Y(\U3/U73/Z_19 ) );
  INVX1 U13283 ( .A(N2899), .Y(n13940) );
  NOR2X1 U13284 ( .A(n12485), .B(n13941), .Y(\U3/U73/Z_18 ) );
  INVX1 U13285 ( .A(N2898), .Y(n13941) );
  NOR2X1 U13286 ( .A(n12485), .B(n13942), .Y(\U3/U73/Z_17 ) );
  INVX1 U13287 ( .A(N2897), .Y(n13942) );
  NOR2X1 U13288 ( .A(n12485), .B(n13943), .Y(\U3/U73/Z_16 ) );
  INVX1 U13289 ( .A(N2896), .Y(n13943) );
  NOR2X1 U13290 ( .A(n12484), .B(n13944), .Y(\U3/U73/Z_15 ) );
  INVX1 U13291 ( .A(N2895), .Y(n13944) );
  AND2X1 U13292 ( .A(N2840), .B(n12477), .Y(\U3/U72/Z_31 ) );
  AND2X1 U13293 ( .A(N2839), .B(n12477), .Y(\U3/U72/Z_30 ) );
  AND2X1 U13294 ( .A(N2838), .B(n12477), .Y(\U3/U72/Z_29 ) );
  AND2X1 U13295 ( .A(N2837), .B(n12477), .Y(\U3/U72/Z_28 ) );
  AND2X1 U13296 ( .A(N2836), .B(n12477), .Y(\U3/U72/Z_27 ) );
  AND2X1 U13297 ( .A(N2835), .B(n12477), .Y(\U3/U72/Z_26 ) );
  AND2X1 U13298 ( .A(N2834), .B(n12477), .Y(\U3/U72/Z_25 ) );
  AND2X1 U13299 ( .A(N2833), .B(n12477), .Y(\U3/U72/Z_24 ) );
  AND2X1 U13300 ( .A(N2832), .B(n12477), .Y(\U3/U72/Z_23 ) );
  AND2X1 U13301 ( .A(N2831), .B(n12477), .Y(\U3/U72/Z_22 ) );
  AND2X1 U13302 ( .A(N2830), .B(n12477), .Y(\U3/U72/Z_21 ) );
  AND2X1 U13303 ( .A(N2829), .B(n12477), .Y(\U3/U72/Z_20 ) );
  AND2X1 U13304 ( .A(N2828), .B(n12477), .Y(\U3/U72/Z_19 ) );
  AND2X1 U13305 ( .A(N2827), .B(n12477), .Y(\U3/U72/Z_18 ) );
  AND2X1 U13306 ( .A(N2826), .B(n12477), .Y(\U3/U72/Z_17 ) );
  AND2X1 U13307 ( .A(N2825), .B(n12477), .Y(\U3/U72/Z_16 ) );
  AND2X1 U13308 ( .A(N2824), .B(n12477), .Y(\U3/U72/Z_15 ) );
  AND2X1 U13309 ( .A(N2171), .B(n12477), .Y(\U3/U71/Z_31 ) );
  AND2X1 U13310 ( .A(N2170), .B(n12477), .Y(\U3/U71/Z_30 ) );
  AND2X1 U13311 ( .A(N2169), .B(n12477), .Y(\U3/U71/Z_29 ) );
  AND2X1 U13312 ( .A(N2168), .B(n12477), .Y(\U3/U71/Z_28 ) );
  AND2X1 U13313 ( .A(N2167), .B(n12477), .Y(\U3/U71/Z_27 ) );
  AND2X1 U13314 ( .A(N2166), .B(n12477), .Y(\U3/U71/Z_26 ) );
  AND2X1 U13315 ( .A(N2165), .B(n12477), .Y(\U3/U71/Z_25 ) );
  AND2X1 U13316 ( .A(N2164), .B(n12477), .Y(\U3/U71/Z_24 ) );
  AND2X1 U13317 ( .A(N2163), .B(n12477), .Y(\U3/U71/Z_23 ) );
  AND2X1 U13318 ( .A(N2162), .B(n12477), .Y(\U3/U71/Z_22 ) );
  AND2X1 U13319 ( .A(N2161), .B(n12477), .Y(\U3/U71/Z_21 ) );
  AND2X1 U13320 ( .A(N2160), .B(n12477), .Y(\U3/U71/Z_20 ) );
  AND2X1 U13321 ( .A(N2159), .B(n12477), .Y(\U3/U71/Z_19 ) );
  AND2X1 U13322 ( .A(N2158), .B(n12477), .Y(\U3/U71/Z_18 ) );
  AND2X1 U13323 ( .A(N2157), .B(n12477), .Y(\U3/U71/Z_17 ) );
  AND2X1 U13324 ( .A(N2156), .B(n12477), .Y(\U3/U71/Z_16 ) );
  AND2X1 U13325 ( .A(N2155), .B(n12477), .Y(\U3/U71/Z_15 ) );
  NOR2X1 U13326 ( .A(n12485), .B(n12755), .Y(\U3/U70/Z_8 ) );
  OAI22X1 U13327 ( .A(n12470), .B(n12732), .C(n12480), .D(n12754), .Y(
        \U3/U70/Z_7 ) );
  OAI22X1 U13328 ( .A(n12470), .B(n12731), .C(n12479), .D(n12753), .Y(
        \U3/U70/Z_6 ) );
  OAI22X1 U13329 ( .A(n12470), .B(n12730), .C(n12479), .D(n12752), .Y(
        \U3/U70/Z_5 ) );
  OAI22X1 U13330 ( .A(n12470), .B(n12729), .C(n12478), .D(n12751), .Y(
        \U3/U70/Z_4 ) );
  OAI22X1 U13331 ( .A(n12470), .B(n12728), .C(n12479), .D(n12750), .Y(
        \U3/U70/Z_3 ) );
  OAI22X1 U13332 ( .A(n12470), .B(n12727), .C(n12478), .D(n12749), .Y(
        \U3/U70/Z_2 ) );
  OAI22X1 U13333 ( .A(n12470), .B(n12726), .C(n12478), .D(n12747), .Y(
        \U3/U70/Z_1 ) );
  NOR2X1 U13334 ( .A(n12470), .B(n12724), .Y(\U3/U70/Z_0 ) );
  AND2X1 U13335 ( .A(N1352), .B(n15370), .Y(\U3/U69/Z_9 ) );
  AND2X1 U13336 ( .A(N1351), .B(n15370), .Y(\U3/U69/Z_8 ) );
  OAI21X1 U13337 ( .A(n12480), .B(n12709), .C(n14328), .Y(\U3/U69/Z_7 ) );
  NAND2X1 U13338 ( .A(N1350), .B(n15370), .Y(n14328) );
  OAI21X1 U13339 ( .A(n12482), .B(n12708), .C(n14329), .Y(\U3/U69/Z_6 ) );
  NAND2X1 U13340 ( .A(N1349), .B(n15370), .Y(n14329) );
  OAI21X1 U13341 ( .A(n12482), .B(n12707), .C(n14330), .Y(\U3/U69/Z_5 ) );
  NAND2X1 U13342 ( .A(N1348), .B(n15370), .Y(n14330) );
  OAI21X1 U13343 ( .A(n12481), .B(n12706), .C(n14331), .Y(\U3/U69/Z_4 ) );
  NAND2X1 U13344 ( .A(N1347), .B(n15370), .Y(n14331) );
  OAI21X1 U13345 ( .A(n12482), .B(n12705), .C(n14332), .Y(\U3/U69/Z_3 ) );
  NAND2X1 U13346 ( .A(N1346), .B(n15370), .Y(n14332) );
  OAI21X1 U13347 ( .A(n12481), .B(n12704), .C(n14333), .Y(\U3/U69/Z_2 ) );
  NAND2X1 U13348 ( .A(N1345), .B(n15370), .Y(n14333) );
  AND2X1 U13349 ( .A(N1356), .B(n15370), .Y(\U3/U69/Z_13 ) );
  AND2X1 U13350 ( .A(N1355), .B(n15370), .Y(\U3/U69/Z_12 ) );
  AND2X1 U13351 ( .A(N1354), .B(n15370), .Y(\U3/U69/Z_11 ) );
  AND2X1 U13352 ( .A(N1353), .B(n15370), .Y(\U3/U69/Z_10 ) );
  OAI21X1 U13353 ( .A(n12481), .B(n12703), .C(n14334), .Y(\U3/U69/Z_1 ) );
  NAND2X1 U13354 ( .A(N1344), .B(n15370), .Y(n14334) );
  OAI21X1 U13355 ( .A(n12482), .B(n12701), .C(n14335), .Y(\U3/U69/Z_0 ) );
  NAND2X1 U13356 ( .A(N1343), .B(n15370), .Y(n14335) );
  AND2X1 U13357 ( .A(N2107), .B(n12477), .Y(\U3/U68/Z_31 ) );
  AND2X1 U13358 ( .A(N2106), .B(n12477), .Y(\U3/U68/Z_30 ) );
  AND2X1 U13359 ( .A(N2105), .B(n12477), .Y(\U3/U68/Z_29 ) );
  AND2X1 U13360 ( .A(N2104), .B(n12477), .Y(\U3/U68/Z_28 ) );
  AND2X1 U13361 ( .A(N2103), .B(n12477), .Y(\U3/U68/Z_27 ) );
  AND2X1 U13362 ( .A(N2102), .B(n12477), .Y(\U3/U68/Z_26 ) );
  AND2X1 U13363 ( .A(N2101), .B(n12477), .Y(\U3/U68/Z_25 ) );
  AND2X1 U13364 ( .A(N2100), .B(n12477), .Y(\U3/U68/Z_24 ) );
  AND2X1 U13365 ( .A(N2099), .B(n12477), .Y(\U3/U68/Z_23 ) );
  AND2X1 U13366 ( .A(N2098), .B(n12477), .Y(\U3/U68/Z_22 ) );
  AND2X1 U13367 ( .A(N2097), .B(n12477), .Y(\U3/U68/Z_21 ) );
  AND2X1 U13368 ( .A(N2096), .B(n12477), .Y(\U3/U68/Z_20 ) );
  AND2X1 U13369 ( .A(N2095), .B(n12477), .Y(\U3/U68/Z_19 ) );
  AND2X1 U13370 ( .A(N2094), .B(n12477), .Y(\U3/U68/Z_18 ) );
  AND2X1 U13371 ( .A(N2093), .B(n12477), .Y(\U3/U68/Z_17 ) );
  AND2X1 U13372 ( .A(N2092), .B(n12477), .Y(\U3/U68/Z_16 ) );
  AND2X1 U13373 ( .A(N2091), .B(n12477), .Y(\U3/U68/Z_15 ) );
  NAND2X1 U13374 ( .A(n12470), .B(n12489), .Y(\U3/U67/Z_1 ) );
  OAI21X1 U13375 ( .A(n12470), .B(n12812), .C(n12486), .Y(\U3/U65/Z_7 ) );
  OAI21X1 U13376 ( .A(n12470), .B(n12811), .C(n12487), .Y(\U3/U65/Z_6 ) );
  OAI21X1 U13377 ( .A(n12470), .B(n12810), .C(n12486), .Y(\U3/U65/Z_5 ) );
  OAI21X1 U13378 ( .A(n12470), .B(n12809), .C(n12486), .Y(\U3/U65/Z_4 ) );
  OAI21X1 U13379 ( .A(n12470), .B(n12808), .C(n12486), .Y(\U3/U65/Z_3 ) );
  OAI21X1 U13380 ( .A(n12470), .B(n12807), .C(n12489), .Y(\U3/U65/Z_2 ) );
  OAI21X1 U13381 ( .A(n12470), .B(n12806), .C(n12489), .Y(\U3/U65/Z_1 ) );
  OAI21X1 U13382 ( .A(n12470), .B(n12804), .C(n12489), .Y(\U3/U65/Z_0 ) );
  NOR2X1 U13383 ( .A(n12486), .B(n12889), .Y(\U3/U64/Z_7 ) );
  NOR2X1 U13384 ( .A(n12485), .B(n12888), .Y(\U3/U64/Z_6 ) );
  NOR2X1 U13385 ( .A(n12486), .B(n12887), .Y(\U3/U64/Z_5 ) );
  NOR2X1 U13386 ( .A(n12486), .B(n12886), .Y(\U3/U64/Z_4 ) );
  NOR2X1 U13387 ( .A(n12486), .B(n12885), .Y(\U3/U64/Z_3 ) );
  NOR2X1 U13388 ( .A(n12485), .B(n12884), .Y(\U3/U64/Z_2 ) );
  NOR2X1 U13389 ( .A(n12478), .B(n12883), .Y(\U3/U64/Z_1 ) );
  OAI21X1 U13390 ( .A(n12480), .B(n12881), .C(n12470), .Y(\U3/U64/Z_0 ) );
  NOR2X1 U13391 ( .A(n12556), .B(n13184), .Y(\U3/U63/Z_7 ) );
  NOR2X1 U13392 ( .A(n12556), .B(n13183), .Y(\U3/U63/Z_6 ) );
  NOR2X1 U13393 ( .A(n12556), .B(n13182), .Y(\U3/U63/Z_5 ) );
  NOR2X1 U13394 ( .A(n12556), .B(n13181), .Y(\U3/U63/Z_4 ) );
  NOR2X1 U13395 ( .A(n12556), .B(n13180), .Y(\U3/U63/Z_3 ) );
  NAND2X1 U13396 ( .A(bCE), .B(n13179), .Y(\U3/U63/Z_2 ) );
  NOR2X1 U13397 ( .A(n12556), .B(n13178), .Y(\U3/U63/Z_1 ) );
  NAND2X1 U13398 ( .A(bCE), .B(n13176), .Y(\U3/U63/Z_0 ) );
  INVX1 U13399 ( .A(n13213), .Y(\U3/U136/Z_0 ) );
  NOR2X1 U13400 ( .A(n12687), .B(n13058), .Y(n13213) );
  NOR2X1 U13401 ( .A(n13905), .B(n12922), .Y(\U3/U134/Z_9 ) );
  INVX1 U13402 ( .A(Gy[9]), .Y(n12922) );
  NOR2X1 U13403 ( .A(n13905), .B(n12920), .Y(\U3/U134/Z_8 ) );
  INVX1 U13404 ( .A(Gy[8]), .Y(n12920) );
  NOR2X1 U13405 ( .A(n13905), .B(n12918), .Y(\U3/U134/Z_7 ) );
  INVX1 U13406 ( .A(Gy[7]), .Y(n12918) );
  NOR2X1 U13407 ( .A(n13905), .B(n12916), .Y(\U3/U134/Z_6 ) );
  INVX1 U13408 ( .A(Gy[6]), .Y(n12916) );
  NOR2X1 U13409 ( .A(n13905), .B(n12914), .Y(\U3/U134/Z_5 ) );
  INVX1 U13410 ( .A(Gy[5]), .Y(n12914) );
  NOR2X1 U13411 ( .A(n13905), .B(n12912), .Y(\U3/U134/Z_4 ) );
  INVX1 U13412 ( .A(Gy[4]), .Y(n12912) );
  NOR2X1 U13413 ( .A(n13905), .B(n12910), .Y(\U3/U134/Z_3 ) );
  INVX1 U13414 ( .A(Gy[3]), .Y(n12910) );
  NOR2X1 U13415 ( .A(n13905), .B(n12908), .Y(\U3/U134/Z_2 ) );
  INVX1 U13416 ( .A(Gy[2]), .Y(n12908) );
  NOR2X1 U13417 ( .A(n13905), .B(n12924), .Y(\U3/U134/Z_10 ) );
  INVX1 U13418 ( .A(Gy[10]), .Y(n12924) );
  NOR2X1 U13419 ( .A(n13905), .B(n12906), .Y(\U3/U134/Z_1 ) );
  INVX1 U13420 ( .A(Gy[1]), .Y(n12906) );
  NOR2X1 U13421 ( .A(n13905), .B(n12903), .Y(\U3/U134/Z_0 ) );
  INVX1 U13422 ( .A(Gy[0]), .Y(n12903) );
  NOR2X1 U13423 ( .A(N2549), .B(n13165), .Y(n13905) );
  OAI21X1 U13424 ( .A(n12470), .B(n12720), .C(n14336), .Y(\U3/U125/Z_7 ) );
  OAI21X1 U13425 ( .A(n12470), .B(n12719), .C(n14336), .Y(\U3/U125/Z_6 ) );
  OAI21X1 U13426 ( .A(n12470), .B(n12718), .C(n14336), .Y(\U3/U125/Z_5 ) );
  OAI21X1 U13427 ( .A(n12470), .B(n12717), .C(n14336), .Y(\U3/U125/Z_4 ) );
  OAI21X1 U13428 ( .A(n12470), .B(n12716), .C(n14336), .Y(\U3/U125/Z_3 ) );
  OAI21X1 U13429 ( .A(n12470), .B(n12715), .C(n14336), .Y(\U3/U125/Z_2 ) );
  OAI21X1 U13430 ( .A(n12470), .B(n12714), .C(n14336), .Y(\U3/U125/Z_1 ) );
  NAND2X1 U13431 ( .A(dy[1]), .B(n15325), .Y(n14336) );
  OAI22X1 U13432 ( .A(n12553), .B(n13419), .C(n12470), .D(n12712), .Y(
        \U3/U125/Z_0 ) );
  INVX1 U13433 ( .A(dy[0]), .Y(n12553) );
  NAND2X1 U13434 ( .A(n13419), .B(n12470), .Y(\U3/U124/Z_0 ) );
  NOR2X1 U13435 ( .A(n13079), .B(n12464), .Y(\U3/U122/Z_9 ) );
  INVX1 U13436 ( .A(fGx[10]), .Y(n13079) );
  NOR2X1 U13437 ( .A(n13063), .B(n13920), .Y(\U3/U122/Z_8 ) );
  INVX1 U13438 ( .A(fGx[9]), .Y(n13063) );
  OAI21X1 U13439 ( .A(n13920), .B(n12970), .C(n14337), .Y(\U3/U122/Z_7 ) );
  OAI21X1 U13440 ( .A(n14338), .B(n14339), .C(n15328), .Y(n14337) );
  NAND2X1 U13441 ( .A(n14340), .B(n14341), .Y(n14339) );
  NOR2X1 U13442 ( .A(n14342), .B(n14343), .Y(n14341) );
  OAI21X1 U13443 ( .A(n12603), .B(n14344), .C(n14345), .Y(n14343) );
  AOI22X1 U13444 ( .A(n14346), .B(N1382), .C(n14347), .D(N1440), .Y(n14345) );
  OAI21X1 U13445 ( .A(n12744), .B(n14348), .C(n14349), .Y(n14342) );
  AOI22X1 U13446 ( .A(n14350), .B(\regX[3][7] ), .C(n14351), .D(\regX[13][7] ), 
        .Y(n14349) );
  INVX1 U13447 ( .A(\regX[5][7] ), .Y(n12744) );
  NOR2X1 U13448 ( .A(n14352), .B(n14353), .Y(n14340) );
  OAI21X1 U13449 ( .A(n12779), .B(n14354), .C(n14355), .Y(n14353) );
  AOI22X1 U13450 ( .A(n14356), .B(\regX[1][7] ), .C(n14357), .D(\regX[11][7] ), 
        .Y(n14355) );
  OAI21X1 U13451 ( .A(n12755), .B(n14358), .C(n14359), .Y(n14352) );
  AOI22X1 U13452 ( .A(n14360), .B(\regX[8][7] ), .C(n14361), .D(N1622), .Y(
        n14359) );
  NAND2X1 U13453 ( .A(n14362), .B(n14363), .Y(n14338) );
  NOR2X1 U13454 ( .A(n14364), .B(n14365), .Y(n14363) );
  OAI21X1 U13455 ( .A(n12860), .B(n14366), .C(n14367), .Y(n14365) );
  AOI22X1 U13456 ( .A(n14368), .B(\regX[16][7] ), .C(n14369), .D(N1742), .Y(
        n14367) );
  OAI21X1 U13457 ( .A(n12801), .B(n14370), .C(n14371), .Y(n14364) );
  AOI22X1 U13458 ( .A(n14372), .B(\regX[22][7] ), .C(n14373), .D(\regX[15][7] ), .Y(n14371) );
  NOR2X1 U13459 ( .A(n14374), .B(n14375), .Y(n14362) );
  OAI21X1 U13460 ( .A(n12850), .B(n14376), .C(n14377), .Y(n14375) );
  AOI22X1 U13461 ( .A(n14378), .B(\regX[24][7] ), .C(n14379), .D(\regX[21][7] ), .Y(n14377) );
  OAI21X1 U13462 ( .A(n13184), .B(n14380), .C(n14381), .Y(n14374) );
  AOI22X1 U13463 ( .A(n14382), .B(\regX[20][7] ), .C(n14383), .D(\regX[18][7] ), .Y(n14381) );
  INVX1 U13464 ( .A(\regX[19][7] ), .Y(n13184) );
  INVX1 U13465 ( .A(fGx[8]), .Y(n12970) );
  OAI21X1 U13466 ( .A(n12464), .B(n14215), .C(n14384), .Y(\U3/U122/Z_6 ) );
  OAI21X1 U13467 ( .A(n14385), .B(n14386), .C(n15328), .Y(n14384) );
  NAND2X1 U13468 ( .A(n14387), .B(n14388), .Y(n14386) );
  NOR2X1 U13469 ( .A(n14389), .B(n14390), .Y(n14388) );
  OAI21X1 U13470 ( .A(n12602), .B(n14344), .C(n14391), .Y(n14390) );
  AOI22X1 U13471 ( .A(n14346), .B(N1381), .C(n14347), .D(N1439), .Y(n14391) );
  OAI21X1 U13472 ( .A(n12743), .B(n14348), .C(n14392), .Y(n14389) );
  AOI22X1 U13473 ( .A(n14350), .B(\regX[3][6] ), .C(n14351), .D(\regX[13][6] ), 
        .Y(n14392) );
  INVX1 U13474 ( .A(\regX[5][6] ), .Y(n12743) );
  NOR2X1 U13475 ( .A(n14393), .B(n14394), .Y(n14387) );
  OAI21X1 U13476 ( .A(n12778), .B(n14354), .C(n14395), .Y(n14394) );
  AOI22X1 U13477 ( .A(n14356), .B(\regX[1][6] ), .C(n14357), .D(\regX[11][6] ), 
        .Y(n14395) );
  OAI21X1 U13478 ( .A(n12754), .B(n14358), .C(n14396), .Y(n14393) );
  AOI22X1 U13479 ( .A(n14360), .B(\regX[8][6] ), .C(n14361), .D(N1621), .Y(
        n14396) );
  NAND2X1 U13480 ( .A(n14397), .B(n14398), .Y(n14385) );
  NOR2X1 U13481 ( .A(n14399), .B(n14400), .Y(n14398) );
  OAI21X1 U13482 ( .A(n12859), .B(n14366), .C(n14401), .Y(n14400) );
  AOI22X1 U13483 ( .A(n14368), .B(\regX[16][6] ), .C(n14369), .D(N1741), .Y(
        n14401) );
  OAI21X1 U13484 ( .A(n12800), .B(n14370), .C(n14402), .Y(n14399) );
  AOI22X1 U13485 ( .A(n14372), .B(\regX[22][6] ), .C(n14373), .D(\regX[15][6] ), .Y(n14402) );
  NOR2X1 U13486 ( .A(n14403), .B(n14404), .Y(n14397) );
  OAI21X1 U13487 ( .A(n12849), .B(n14376), .C(n14405), .Y(n14404) );
  AOI22X1 U13488 ( .A(n14378), .B(\regX[24][6] ), .C(n14379), .D(\regX[21][6] ), .Y(n14405) );
  OAI21X1 U13489 ( .A(n13183), .B(n14380), .C(n14406), .Y(n14403) );
  AOI22X1 U13490 ( .A(n14382), .B(\regX[20][6] ), .C(n14383), .D(\regX[18][6] ), .Y(n14406) );
  INVX1 U13491 ( .A(\regX[19][6] ), .Y(n13183) );
  INVX1 U13492 ( .A(fGx[7]), .Y(n14215) );
  OAI21X1 U13493 ( .A(n13920), .B(n14217), .C(n14407), .Y(\U3/U122/Z_5 ) );
  OAI21X1 U13494 ( .A(n14408), .B(n14409), .C(n15328), .Y(n14407) );
  NAND2X1 U13495 ( .A(n14410), .B(n14411), .Y(n14409) );
  NOR2X1 U13496 ( .A(n14412), .B(n14413), .Y(n14411) );
  OAI21X1 U13497 ( .A(n12601), .B(n14344), .C(n14414), .Y(n14413) );
  AOI22X1 U13498 ( .A(n14346), .B(N1380), .C(n14347), .D(N1438), .Y(n14414) );
  OAI21X1 U13499 ( .A(n12742), .B(n14348), .C(n14415), .Y(n14412) );
  AOI22X1 U13500 ( .A(n14350), .B(\regX[3][5] ), .C(n14351), .D(\regX[13][5] ), 
        .Y(n14415) );
  INVX1 U13501 ( .A(\regX[5][5] ), .Y(n12742) );
  NOR2X1 U13502 ( .A(n14416), .B(n14417), .Y(n14410) );
  OAI21X1 U13503 ( .A(n12777), .B(n14354), .C(n14418), .Y(n14417) );
  AOI22X1 U13504 ( .A(n14356), .B(\regX[1][5] ), .C(n14357), .D(\regX[11][5] ), 
        .Y(n14418) );
  OAI21X1 U13505 ( .A(n12753), .B(n14358), .C(n14419), .Y(n14416) );
  AOI22X1 U13506 ( .A(n14360), .B(\regX[8][5] ), .C(n14361), .D(N1620), .Y(
        n14419) );
  NAND2X1 U13507 ( .A(n14420), .B(n14421), .Y(n14408) );
  NOR2X1 U13508 ( .A(n14422), .B(n14423), .Y(n14421) );
  OAI21X1 U13509 ( .A(n12858), .B(n14366), .C(n14424), .Y(n14423) );
  AOI22X1 U13510 ( .A(n14368), .B(\regX[16][5] ), .C(n14369), .D(N1740), .Y(
        n14424) );
  OAI21X1 U13511 ( .A(n12799), .B(n14370), .C(n14425), .Y(n14422) );
  AOI22X1 U13512 ( .A(n14372), .B(\regX[22][5] ), .C(n14373), .D(\regX[15][5] ), .Y(n14425) );
  NOR2X1 U13513 ( .A(n14426), .B(n14427), .Y(n14420) );
  OAI21X1 U13514 ( .A(n12848), .B(n14376), .C(n14428), .Y(n14427) );
  AOI22X1 U13515 ( .A(n14378), .B(\regX[24][5] ), .C(n14379), .D(\regX[21][5] ), .Y(n14428) );
  OAI21X1 U13516 ( .A(n13182), .B(n14380), .C(n14429), .Y(n14426) );
  AOI22X1 U13517 ( .A(n14382), .B(\regX[20][5] ), .C(n14383), .D(\regX[18][5] ), .Y(n14429) );
  INVX1 U13518 ( .A(\regX[19][5] ), .Y(n13182) );
  INVX1 U13519 ( .A(fGx[6]), .Y(n14217) );
  OAI21X1 U13520 ( .A(n12464), .B(n14219), .C(n14430), .Y(\U3/U122/Z_4 ) );
  OAI21X1 U13521 ( .A(n14431), .B(n14432), .C(n15328), .Y(n14430) );
  NAND2X1 U13522 ( .A(n14433), .B(n14434), .Y(n14432) );
  NOR2X1 U13523 ( .A(n14435), .B(n14436), .Y(n14434) );
  OAI21X1 U13524 ( .A(n12600), .B(n14344), .C(n14437), .Y(n14436) );
  AOI22X1 U13525 ( .A(n14346), .B(N1379), .C(n14347), .D(N1437), .Y(n14437) );
  INVX1 U13526 ( .A(n14438), .Y(n14347) );
  OAI21X1 U13527 ( .A(n12741), .B(n14348), .C(n14439), .Y(n14435) );
  AOI22X1 U13528 ( .A(n14350), .B(\regX[3][4] ), .C(n14351), .D(\regX[13][4] ), 
        .Y(n14439) );
  INVX1 U13529 ( .A(n14440), .Y(n14350) );
  INVX1 U13530 ( .A(\regX[5][4] ), .Y(n12741) );
  NOR2X1 U13531 ( .A(n14441), .B(n14442), .Y(n14433) );
  OAI21X1 U13532 ( .A(n12776), .B(n14354), .C(n14443), .Y(n14442) );
  AOI22X1 U13533 ( .A(n14356), .B(\regX[1][4] ), .C(n14357), .D(\regX[11][4] ), 
        .Y(n14443) );
  OAI21X1 U13534 ( .A(n12752), .B(n14358), .C(n14444), .Y(n14441) );
  AOI22X1 U13535 ( .A(n14360), .B(\regX[8][4] ), .C(n14361), .D(N1619), .Y(
        n14444) );
  NAND2X1 U13536 ( .A(n14445), .B(n14446), .Y(n14431) );
  NOR2X1 U13537 ( .A(n14447), .B(n14448), .Y(n14446) );
  OAI21X1 U13538 ( .A(n12857), .B(n14366), .C(n14449), .Y(n14448) );
  AOI22X1 U13539 ( .A(n14368), .B(\regX[16][4] ), .C(n14369), .D(N1739), .Y(
        n14449) );
  OAI21X1 U13540 ( .A(n12798), .B(n14370), .C(n14450), .Y(n14447) );
  AOI22X1 U13541 ( .A(n14372), .B(\regX[22][4] ), .C(n14373), .D(\regX[15][4] ), .Y(n14450) );
  INVX1 U13542 ( .A(n14451), .Y(n14372) );
  NOR2X1 U13543 ( .A(n14452), .B(n14453), .Y(n14445) );
  OAI21X1 U13544 ( .A(n12847), .B(n14376), .C(n14454), .Y(n14453) );
  AOI22X1 U13545 ( .A(n14378), .B(\regX[24][4] ), .C(n14379), .D(\regX[21][4] ), .Y(n14454) );
  INVX1 U13546 ( .A(n14455), .Y(n14379) );
  OAI21X1 U13547 ( .A(n13181), .B(n14380), .C(n14456), .Y(n14452) );
  AOI22X1 U13548 ( .A(n14382), .B(\regX[20][4] ), .C(n14383), .D(\regX[18][4] ), .Y(n14456) );
  INVX1 U13549 ( .A(n14457), .Y(n14382) );
  INVX1 U13550 ( .A(\regX[19][4] ), .Y(n13181) );
  INVX1 U13551 ( .A(fGx[5]), .Y(n14219) );
  OAI21X1 U13552 ( .A(n13920), .B(n14221), .C(n14458), .Y(\U3/U122/Z_3 ) );
  OAI21X1 U13553 ( .A(n14459), .B(n14460), .C(n15328), .Y(n14458) );
  NAND2X1 U13554 ( .A(n14461), .B(n14462), .Y(n14460) );
  NOR2X1 U13555 ( .A(n14463), .B(n14464), .Y(n14462) );
  OAI21X1 U13556 ( .A(n12751), .B(n14358), .C(n14465), .Y(n14464) );
  AOI22X1 U13557 ( .A(n14356), .B(\regX[1][3] ), .C(n14357), .D(\regX[11][3] ), 
        .Y(n14465) );
  INVX1 U13558 ( .A(\regX[7][3] ), .Y(n12751) );
  OAI21X1 U13559 ( .A(n12846), .B(n14376), .C(n14466), .Y(n14463) );
  AOI22X1 U13560 ( .A(n14360), .B(\regX[8][3] ), .C(n14361), .D(N1618), .Y(
        n14466) );
  NOR2X1 U13561 ( .A(n14467), .B(n14468), .Y(n14461) );
  OAI21X1 U13562 ( .A(n12775), .B(n14354), .C(n14469), .Y(n14468) );
  AOI22X1 U13563 ( .A(n14470), .B(\regX[5][3] ), .C(n14471), .D(\regX[0][3] ), 
        .Y(n14469) );
  OAI21X1 U13564 ( .A(n12728), .B(n14438), .C(n14472), .Y(n14467) );
  AOI22X1 U13565 ( .A(n14346), .B(N1378), .C(n14351), .D(\regX[13][3] ), .Y(
        n14472) );
  INVX1 U13566 ( .A(N1436), .Y(n12728) );
  NAND3X1 U13567 ( .A(n14473), .B(n14474), .C(n14475), .Y(n14459) );
  NOR2X1 U13568 ( .A(n14476), .B(n14477), .Y(n14475) );
  OAI21X1 U13569 ( .A(n12797), .B(n14370), .C(n14478), .Y(n14477) );
  AOI22X1 U13570 ( .A(n14373), .B(\regX[15][3] ), .C(n14479), .D(N1680), .Y(
        n14478) );
  INVX1 U13571 ( .A(\regX[17][3] ), .Y(n12797) );
  OAI21X1 U13572 ( .A(n13180), .B(n14380), .C(n14480), .Y(n14476) );
  AOI22X1 U13573 ( .A(n14368), .B(\regX[16][3] ), .C(n14369), .D(N1738), .Y(
        n14480) );
  INVX1 U13574 ( .A(\regX[19][3] ), .Y(n13180) );
  NOR2X1 U13575 ( .A(n14481), .B(n14482), .Y(n14474) );
  OAI22X1 U13576 ( .A(n12836), .B(n14451), .C(n12865), .D(n14457), .Y(n14482)
         );
  INVX1 U13577 ( .A(\regX[20][3] ), .Y(n12865) );
  INVX1 U13578 ( .A(\regX[22][3] ), .Y(n12836) );
  OAI22X1 U13579 ( .A(n12808), .B(n14483), .C(n12673), .D(n14484), .Y(n14481)
         );
  INVX1 U13580 ( .A(\regX[24][3] ), .Y(n12808) );
  AOI21X1 U13581 ( .A(n14383), .B(\regX[18][3] ), .C(n14485), .Y(n14473) );
  OAI22X1 U13582 ( .A(n12875), .B(n14455), .C(n12716), .D(n14440), .Y(n14485)
         );
  INVX1 U13583 ( .A(\regX[3][3] ), .Y(n12716) );
  INVX1 U13584 ( .A(fGx[4]), .Y(n14221) );
  NOR2X1 U13585 ( .A(n13159), .B(n12464), .Y(\U3/U122/Z_29 ) );
  INVX1 U13586 ( .A(fGx[30]), .Y(n13159) );
  NOR2X1 U13587 ( .A(n13155), .B(n13920), .Y(\U3/U122/Z_28 ) );
  INVX1 U13588 ( .A(fGx[29]), .Y(n13155) );
  NOR2X1 U13589 ( .A(n13151), .B(n12464), .Y(\U3/U122/Z_27 ) );
  INVX1 U13590 ( .A(fGx[28]), .Y(n13151) );
  NOR2X1 U13591 ( .A(n13147), .B(n13920), .Y(\U3/U122/Z_26 ) );
  INVX1 U13592 ( .A(fGx[27]), .Y(n13147) );
  NOR2X1 U13593 ( .A(n13143), .B(n12464), .Y(\U3/U122/Z_25 ) );
  INVX1 U13594 ( .A(fGx[26]), .Y(n13143) );
  NOR2X1 U13595 ( .A(n13139), .B(n13920), .Y(\U3/U122/Z_24 ) );
  INVX1 U13596 ( .A(fGx[25]), .Y(n13139) );
  NOR2X1 U13597 ( .A(n13135), .B(n12464), .Y(\U3/U122/Z_23 ) );
  INVX1 U13598 ( .A(fGx[24]), .Y(n13135) );
  NOR2X1 U13599 ( .A(n13131), .B(n13920), .Y(\U3/U122/Z_22 ) );
  INVX1 U13600 ( .A(fGx[23]), .Y(n13131) );
  NOR2X1 U13601 ( .A(n13127), .B(n12464), .Y(\U3/U122/Z_21 ) );
  INVX1 U13602 ( .A(fGx[22]), .Y(n13127) );
  NOR2X1 U13603 ( .A(n13123), .B(n13920), .Y(\U3/U122/Z_20 ) );
  INVX1 U13604 ( .A(fGx[21]), .Y(n13123) );
  OAI21X1 U13605 ( .A(n12464), .B(n14223), .C(n14486), .Y(\U3/U122/Z_2 ) );
  OAI21X1 U13606 ( .A(n14487), .B(n14488), .C(n15328), .Y(n14486) );
  NAND2X1 U13607 ( .A(n14489), .B(n14490), .Y(n14488) );
  NOR2X1 U13608 ( .A(n14491), .B(n14492), .Y(n14490) );
  OAI21X1 U13609 ( .A(n12750), .B(n14358), .C(n14493), .Y(n14492) );
  AOI22X1 U13610 ( .A(n14356), .B(\regX[1][2] ), .C(n14357), .D(\regX[11][2] ), 
        .Y(n14493) );
  INVX1 U13611 ( .A(\regX[7][2] ), .Y(n12750) );
  OAI21X1 U13612 ( .A(n12845), .B(n14376), .C(n14494), .Y(n14491) );
  AOI22X1 U13613 ( .A(n14360), .B(\regX[8][2] ), .C(n14361), .D(N1617), .Y(
        n14494) );
  NOR2X1 U13614 ( .A(n14495), .B(n14496), .Y(n14489) );
  OAI21X1 U13615 ( .A(n12774), .B(n14354), .C(n14497), .Y(n14496) );
  AOI22X1 U13616 ( .A(n14470), .B(\regX[5][2] ), .C(n14471), .D(\regX[0][2] ), 
        .Y(n14497) );
  OAI21X1 U13617 ( .A(n12727), .B(n14438), .C(n14498), .Y(n14495) );
  AOI22X1 U13618 ( .A(n14346), .B(N1377), .C(n14351), .D(\regX[13][2] ), .Y(
        n14498) );
  INVX1 U13619 ( .A(N1435), .Y(n12727) );
  NAND3X1 U13620 ( .A(n14499), .B(n14500), .C(n14501), .Y(n14487) );
  NOR2X1 U13621 ( .A(n14502), .B(n14503), .Y(n14501) );
  OAI21X1 U13622 ( .A(n12796), .B(n14370), .C(n14504), .Y(n14503) );
  AOI22X1 U13623 ( .A(n14373), .B(\regX[15][2] ), .C(n14479), .D(N1679), .Y(
        n14504) );
  INVX1 U13624 ( .A(\regX[17][2] ), .Y(n12796) );
  OAI21X1 U13625 ( .A(n13179), .B(n14380), .C(n14505), .Y(n14502) );
  AOI22X1 U13626 ( .A(n14368), .B(\regX[16][2] ), .C(n14369), .D(N1737), .Y(
        n14505) );
  INVX1 U13627 ( .A(\regX[19][2] ), .Y(n13179) );
  NOR2X1 U13628 ( .A(n14506), .B(n14507), .Y(n14500) );
  OAI22X1 U13629 ( .A(n12835), .B(n14451), .C(n12864), .D(n14457), .Y(n14507)
         );
  OAI22X1 U13630 ( .A(n12807), .B(n14483), .C(n12672), .D(n14484), .Y(n14506)
         );
  AOI21X1 U13631 ( .A(n14383), .B(\regX[18][2] ), .C(n14508), .Y(n14499) );
  OAI22X1 U13632 ( .A(n12874), .B(n14455), .C(n12715), .D(n14440), .Y(n14508)
         );
  INVX1 U13633 ( .A(fGx[3]), .Y(n14223) );
  NOR2X1 U13634 ( .A(n13119), .B(n12464), .Y(\U3/U122/Z_19 ) );
  INVX1 U13635 ( .A(fGx[20]), .Y(n13119) );
  NOR2X1 U13636 ( .A(n13115), .B(n13920), .Y(\U3/U122/Z_18 ) );
  INVX1 U13637 ( .A(fGx[19]), .Y(n13115) );
  NOR2X1 U13638 ( .A(n13111), .B(n12464), .Y(\U3/U122/Z_17 ) );
  INVX1 U13639 ( .A(fGx[18]), .Y(n13111) );
  NOR2X1 U13640 ( .A(n13107), .B(n13920), .Y(\U3/U122/Z_16 ) );
  INVX1 U13641 ( .A(fGx[17]), .Y(n13107) );
  NOR2X1 U13642 ( .A(n13103), .B(n12464), .Y(\U3/U122/Z_15 ) );
  INVX1 U13643 ( .A(fGx[16]), .Y(n13103) );
  NOR2X1 U13644 ( .A(n13099), .B(n13920), .Y(\U3/U122/Z_14 ) );
  INVX1 U13645 ( .A(fGx[15]), .Y(n13099) );
  NOR2X1 U13646 ( .A(n13095), .B(n12464), .Y(\U3/U122/Z_13 ) );
  INVX1 U13647 ( .A(fGx[14]), .Y(n13095) );
  NOR2X1 U13648 ( .A(n13091), .B(n13920), .Y(\U3/U122/Z_12 ) );
  INVX1 U13649 ( .A(fGx[13]), .Y(n13091) );
  NOR2X1 U13650 ( .A(n13087), .B(n12464), .Y(\U3/U122/Z_11 ) );
  INVX1 U13651 ( .A(fGx[12]), .Y(n13087) );
  NOR2X1 U13652 ( .A(n13083), .B(n13920), .Y(\U3/U122/Z_10 ) );
  INVX1 U13653 ( .A(fGx[11]), .Y(n13083) );
  OAI21X1 U13654 ( .A(n13920), .B(n14225), .C(n14509), .Y(\U3/U122/Z_1 ) );
  OAI21X1 U13655 ( .A(n14510), .B(n14511), .C(n15328), .Y(n14509) );
  NAND2X1 U13656 ( .A(n14512), .B(n14513), .Y(n14511) );
  NOR2X1 U13657 ( .A(n14514), .B(n14515), .Y(n14513) );
  OAI21X1 U13658 ( .A(n12749), .B(n14358), .C(n14516), .Y(n14515) );
  AOI22X1 U13659 ( .A(n14356), .B(\regX[1][1] ), .C(n14357), .D(\regX[11][1] ), 
        .Y(n14516) );
  INVX1 U13660 ( .A(\regX[7][1] ), .Y(n12749) );
  OAI21X1 U13661 ( .A(n12844), .B(n14376), .C(n14517), .Y(n14514) );
  AOI22X1 U13662 ( .A(n14360), .B(\regX[8][1] ), .C(n14361), .D(N1616), .Y(
        n14517) );
  NOR2X1 U13663 ( .A(n14518), .B(n14519), .Y(n14512) );
  OAI21X1 U13664 ( .A(n12773), .B(n14354), .C(n14520), .Y(n14519) );
  AOI22X1 U13665 ( .A(n14470), .B(\regX[5][1] ), .C(n14471), .D(\regX[0][1] ), 
        .Y(n14520) );
  OAI21X1 U13666 ( .A(n12726), .B(n14438), .C(n14521), .Y(n14518) );
  AOI22X1 U13667 ( .A(n14346), .B(N1376), .C(n14351), .D(\regX[13][1] ), .Y(
        n14521) );
  INVX1 U13668 ( .A(N1434), .Y(n12726) );
  NAND3X1 U13669 ( .A(n14522), .B(n14523), .C(n14524), .Y(n14510) );
  NOR2X1 U13670 ( .A(n14525), .B(n14526), .Y(n14524) );
  OAI21X1 U13671 ( .A(n12795), .B(n14370), .C(n14527), .Y(n14526) );
  AOI22X1 U13672 ( .A(n14373), .B(\regX[15][1] ), .C(n14479), .D(N1678), .Y(
        n14527) );
  INVX1 U13673 ( .A(\regX[17][1] ), .Y(n12795) );
  OAI21X1 U13674 ( .A(n13178), .B(n14380), .C(n14528), .Y(n14525) );
  AOI22X1 U13675 ( .A(n14368), .B(\regX[16][1] ), .C(n14369), .D(N1736), .Y(
        n14528) );
  INVX1 U13676 ( .A(\regX[19][1] ), .Y(n13178) );
  NOR2X1 U13677 ( .A(n14529), .B(n14530), .Y(n14523) );
  OAI22X1 U13678 ( .A(n12834), .B(n14451), .C(n12863), .D(n14457), .Y(n14530)
         );
  INVX1 U13679 ( .A(\regX[20][1] ), .Y(n12863) );
  INVX1 U13680 ( .A(\regX[22][1] ), .Y(n12834) );
  OAI22X1 U13681 ( .A(n12806), .B(n14483), .C(n12671), .D(n14484), .Y(n14529)
         );
  INVX1 U13682 ( .A(\regX[24][1] ), .Y(n12806) );
  AOI21X1 U13683 ( .A(n14383), .B(\regX[18][1] ), .C(n14531), .Y(n14522) );
  OAI22X1 U13684 ( .A(n12873), .B(n14455), .C(n12714), .D(n14440), .Y(n14531)
         );
  INVX1 U13685 ( .A(\regX[3][1] ), .Y(n12714) );
  INVX1 U13686 ( .A(fGx[2]), .Y(n14225) );
  OAI21X1 U13687 ( .A(n12464), .B(n14227), .C(n14532), .Y(\U3/U122/Z_0 ) );
  OAI21X1 U13688 ( .A(n14533), .B(n14534), .C(n15328), .Y(n14532) );
  NAND2X1 U13689 ( .A(n14535), .B(n14536), .Y(n14534) );
  NOR2X1 U13690 ( .A(n14537), .B(n14538), .Y(n14536) );
  OAI21X1 U13691 ( .A(n12747), .B(n14358), .C(n14539), .Y(n14538) );
  AOI22X1 U13692 ( .A(n14356), .B(\regX[1][0] ), .C(n14357), .D(\regX[11][0] ), 
        .Y(n14539) );
  AND2X1 U13693 ( .A(n14540), .B(n14541), .Y(n14357) );
  AND2X1 U13694 ( .A(n14542), .B(n14543), .Y(n14356) );
  NAND2X1 U13695 ( .A(n14542), .B(n14544), .Y(n14358) );
  INVX1 U13696 ( .A(\regX[7][0] ), .Y(n12747) );
  OAI21X1 U13697 ( .A(n12842), .B(n14376), .C(n14545), .Y(n14537) );
  AOI22X1 U13698 ( .A(n14360), .B(\regX[8][0] ), .C(n14361), .D(N1615), .Y(
        n14545) );
  AND2X1 U13699 ( .A(n14540), .B(n14546), .Y(n14361) );
  INVX1 U13700 ( .A(n14547), .Y(n14360) );
  NAND3X1 U13701 ( .A(n14546), .B(n14543), .C(n14548), .Y(n14547) );
  NAND2X1 U13702 ( .A(n14549), .B(n14544), .Y(n14376) );
  NOR2X1 U13703 ( .A(n14550), .B(n14551), .Y(n14535) );
  OAI21X1 U13704 ( .A(n12771), .B(n14354), .C(n14552), .Y(n14551) );
  AOI22X1 U13705 ( .A(n14470), .B(\regX[5][0] ), .C(n14471), .D(\regX[0][0] ), 
        .Y(n14552) );
  INVX1 U13706 ( .A(n14344), .Y(n14471) );
  NAND2X1 U13707 ( .A(n14553), .B(n14543), .Y(n14344) );
  INVX1 U13708 ( .A(n14348), .Y(n14470) );
  NAND2X1 U13709 ( .A(n14542), .B(n14554), .Y(n14348) );
  NAND2X1 U13710 ( .A(n14543), .B(n14541), .Y(n14354) );
  OAI21X1 U13711 ( .A(n12724), .B(n14438), .C(n14555), .Y(n14550) );
  AOI22X1 U13712 ( .A(n14346), .B(N1375), .C(n14351), .D(\regX[13][0] ), .Y(
        n14555) );
  AND2X1 U13713 ( .A(n14554), .B(n14541), .Y(n14351) );
  AND2X1 U13714 ( .A(n14553), .B(n14540), .Y(n14346) );
  NAND2X1 U13715 ( .A(n14553), .B(n14554), .Y(n14438) );
  INVX1 U13716 ( .A(N1433), .Y(n12724) );
  NAND3X1 U13717 ( .A(n14556), .B(n14557), .C(n14558), .Y(n14533) );
  NOR2X1 U13718 ( .A(n14559), .B(n14560), .Y(n14558) );
  OAI21X1 U13719 ( .A(n12793), .B(n14370), .C(n14561), .Y(n14560) );
  AOI22X1 U13720 ( .A(n14373), .B(\regX[15][0] ), .C(n14479), .D(N1677), .Y(
        n14561) );
  INVX1 U13721 ( .A(n14366), .Y(n14479) );
  NAND2X1 U13722 ( .A(n14554), .B(n14546), .Y(n14366) );
  AND2X1 U13723 ( .A(n14541), .B(n14544), .Y(n14373) );
  NOR2X1 U13724 ( .A(n14562), .B(n14563), .Y(n14541) );
  NAND2X1 U13725 ( .A(n14543), .B(n14549), .Y(n14370) );
  INVX1 U13726 ( .A(\regX[17][0] ), .Y(n12793) );
  OAI21X1 U13727 ( .A(n13176), .B(n14380), .C(n14564), .Y(n14559) );
  AOI22X1 U13728 ( .A(n14368), .B(\regX[16][0] ), .C(n14369), .D(N1735), .Y(
        n14564) );
  AND2X1 U13729 ( .A(n14546), .B(n14544), .Y(n14369) );
  NOR2X1 U13730 ( .A(n14562), .B(n14565), .Y(n14546) );
  INVX1 U13731 ( .A(n14566), .Y(n14368) );
  NAND3X1 U13732 ( .A(n14567), .B(n14562), .C(n14543), .Y(n14566) );
  NOR2X1 U13733 ( .A(n14568), .B(n14569), .Y(n14543) );
  NAND2X1 U13734 ( .A(n14540), .B(n14549), .Y(n14380) );
  INVX1 U13735 ( .A(\regX[19][0] ), .Y(n13176) );
  NOR2X1 U13736 ( .A(n14570), .B(n14571), .Y(n14557) );
  OAI22X1 U13737 ( .A(n12832), .B(n14451), .C(n12861), .D(n14457), .Y(n14571)
         );
  NAND2X1 U13738 ( .A(n14554), .B(n14567), .Y(n14457) );
  NAND2X1 U13739 ( .A(n14544), .B(n14567), .Y(n14451) );
  OAI22X1 U13740 ( .A(n12804), .B(n14483), .C(n12669), .D(n14484), .Y(n14570)
         );
  NAND2X1 U13741 ( .A(n14553), .B(n14544), .Y(n14484) );
  NOR2X1 U13742 ( .A(n14572), .B(n14573), .Y(n14544) );
  INVX1 U13743 ( .A(n14574), .Y(n14553) );
  NAND3X1 U13744 ( .A(n14563), .B(n14562), .C(n14548), .Y(n14574) );
  INVX1 U13745 ( .A(n14378), .Y(n14483) );
  NOR2X1 U13746 ( .A(n14562), .B(n14548), .Y(n14378) );
  AOI21X1 U13747 ( .A(n14383), .B(\regX[18][0] ), .C(n14575), .Y(n14556) );
  OAI22X1 U13748 ( .A(n12871), .B(n14455), .C(n12712), .D(n14440), .Y(n14575)
         );
  NAND2X1 U13749 ( .A(n14542), .B(n14540), .Y(n14440) );
  INVX1 U13750 ( .A(n14576), .Y(n14542) );
  NAND3X1 U13751 ( .A(n14562), .B(n14565), .C(n14548), .Y(n14576) );
  NAND2X1 U13752 ( .A(n14554), .B(n14549), .Y(n14455) );
  NOR2X1 U13753 ( .A(n14563), .B(n14548), .Y(n14549) );
  NOR2X1 U13754 ( .A(n14573), .B(n14569), .Y(n14554) );
  AND2X1 U13755 ( .A(n14540), .B(n14567), .Y(n14383) );
  NOR2X1 U13756 ( .A(n14565), .B(n14548), .Y(n14567) );
  XOR2X1 U13757 ( .A(n14577), .B(n14578), .Y(n14548) );
  XNOR2X1 U13758 ( .A(n14579), .B(n14183), .Y(n14577) );
  XOR2X1 U13759 ( .A(n14580), .B(n14581), .Y(n14183) );
  AOI21X1 U13760 ( .A(n15369), .B(N3093), .C(n14582), .Y(n14581) );
  NAND2X1 U13761 ( .A(n14583), .B(n14584), .Y(n14580) );
  OAI21X1 U13762 ( .A(n14585), .B(n14586), .C(n14587), .Y(n14583) );
  OAI21X1 U13763 ( .A(n14588), .B(n14589), .C(n14590), .Y(n14579) );
  OAI21X1 U13764 ( .A(n14591), .B(n14592), .C(n14578), .Y(n14590) );
  INVX1 U13765 ( .A(n14591), .Y(n14589) );
  NOR2X1 U13766 ( .A(n14572), .B(n14568), .Y(n14540) );
  INVX1 U13767 ( .A(n14573), .Y(n14568) );
  XNOR2X1 U13768 ( .A(n14593), .B(n14578), .Y(n14573) );
  XNOR2X1 U13769 ( .A(n14200), .B(n14594), .Y(n14593) );
  INVX1 U13770 ( .A(fGx[1]), .Y(n14227) );
  AND2X1 U13771 ( .A(fGy[7]), .B(n12466), .Y(\U3/U121/Z_7 ) );
  AND2X1 U13772 ( .A(fGy[6]), .B(n12466), .Y(\U3/U121/Z_6 ) );
  AND2X1 U13773 ( .A(fGy[5]), .B(n12466), .Y(\U3/U121/Z_5 ) );
  AND2X1 U13774 ( .A(fGy[4]), .B(n12466), .Y(\U3/U121/Z_4 ) );
  OAI21X1 U13775 ( .A(n13920), .B(n14595), .C(n12552), .Y(\U3/U121/Z_3 ) );
  OAI21X1 U13776 ( .A(n12464), .B(n14596), .C(n12552), .Y(\U3/U121/Z_2 ) );
  OAI21X1 U13777 ( .A(n13920), .B(n14597), .C(n12552), .Y(\U3/U121/Z_1 ) );
  OAI21X1 U13778 ( .A(n13920), .B(n14598), .C(n12552), .Y(\U3/U121/Z_0 ) );
  INVX1 U13779 ( .A(n12466), .Y(n13920) );
  NOR2X1 U13780 ( .A(n14214), .B(n14318), .Y(\U3/U119/Z_9 ) );
  INVX1 U13781 ( .A(N2755), .Y(n14318) );
  NOR2X1 U13782 ( .A(n14214), .B(n14294), .Y(\U3/U119/Z_8 ) );
  INVX1 U13783 ( .A(N2754), .Y(n14294) );
  NAND3X1 U13784 ( .A(n14599), .B(n14600), .C(n14601), .Y(\U3/U119/Z_7 ) );
  NOR2X1 U13785 ( .A(n14602), .B(n14603), .Y(n14601) );
  OR2X1 U13786 ( .A(n14604), .B(n14605), .Y(n14603) );
  OAI21X1 U13787 ( .A(n12801), .B(n14606), .C(n14607), .Y(n14605) );
  AOI22X1 U13788 ( .A(n14608), .B(\regX[16][7] ), .C(n14609), .D(\regX[24][7] ), .Y(n14607) );
  INVX1 U13789 ( .A(\regX[17][7] ), .Y(n12801) );
  OAI21X1 U13790 ( .A(n12732), .B(n14610), .C(n14611), .Y(n14604) );
  AOI22X1 U13791 ( .A(n14612), .B(\regX[15][7] ), .C(n14613), .D(N1742), .Y(
        n14611) );
  INVX1 U13792 ( .A(N1440), .Y(n12732) );
  NAND3X1 U13793 ( .A(n14614), .B(n14615), .C(n14616), .Y(n14602) );
  AOI21X1 U13794 ( .A(n14617), .B(\regX[21][7] ), .C(n14618), .Y(n14616) );
  OAI22X1 U13795 ( .A(n12850), .B(n14619), .C(n13174), .D(n14620), .Y(n14618)
         );
  INVX1 U13796 ( .A(\regX[23][7] ), .Y(n12850) );
  AOI22X1 U13797 ( .A(n14621), .B(N1684), .C(n14622), .D(\regX[19][7] ), .Y(
        n14615) );
  AOI22X1 U13798 ( .A(n14623), .B(\regX[13][7] ), .C(n14624), .D(\regX[20][7] ), .Y(n14614) );
  NOR2X1 U13799 ( .A(n14625), .B(n14626), .Y(n14600) );
  OAI21X1 U13800 ( .A(n12603), .B(n14627), .C(n14628), .Y(n14626) );
  AOI22X1 U13801 ( .A(n14629), .B(\regX[22][7] ), .C(n14630), .D(\regX[1][7] ), 
        .Y(n14628) );
  INVX1 U13802 ( .A(\regX[0][7] ), .Y(n12603) );
  OR2X1 U13803 ( .A(n14631), .B(n14632), .Y(n14625) );
  OAI22X1 U13804 ( .A(n12768), .B(n14633), .C(n12779), .D(n14634), .Y(n14632)
         );
  OAI21X1 U13805 ( .A(n12755), .B(n14635), .C(n12505), .Y(n14631) );
  NAND2X1 U13806 ( .A(N2753), .B(n15377), .Y(n12505) );
  INVX1 U13807 ( .A(\regX[7][7] ), .Y(n12755) );
  NOR2X1 U13808 ( .A(n14636), .B(n14637), .Y(n14599) );
  OAI21X1 U13809 ( .A(n12720), .B(n14638), .C(n14639), .Y(n14637) );
  AOI22X1 U13810 ( .A(n14640), .B(N1382), .C(\regX[6][7] ), .D(n14641), .Y(
        n14639) );
  OAI21X1 U13811 ( .A(n12899), .B(n14642), .C(n14643), .Y(n14636) );
  AOI22X1 U13812 ( .A(n14644), .B(\regX[5][7] ), .C(n14645), .D(N1622), .Y(
        n14643) );
  INVX1 U13813 ( .A(\regX[11][7] ), .Y(n12899) );
  NAND3X1 U13814 ( .A(n14646), .B(n14647), .C(n14648), .Y(\U3/U119/Z_6 ) );
  NOR2X1 U13815 ( .A(n14649), .B(n14650), .Y(n14648) );
  OR2X1 U13816 ( .A(n14651), .B(n14652), .Y(n14650) );
  OAI21X1 U13817 ( .A(n12800), .B(n14606), .C(n14653), .Y(n14652) );
  AOI22X1 U13818 ( .A(n14608), .B(\regX[16][6] ), .C(n14609), .D(\regX[24][6] ), .Y(n14653) );
  INVX1 U13819 ( .A(\regX[17][6] ), .Y(n12800) );
  OAI21X1 U13820 ( .A(n12731), .B(n14610), .C(n14654), .Y(n14651) );
  AOI22X1 U13821 ( .A(n14612), .B(\regX[15][6] ), .C(n14613), .D(N1741), .Y(
        n14654) );
  INVX1 U13822 ( .A(N1439), .Y(n12731) );
  NAND3X1 U13823 ( .A(n14655), .B(n14656), .C(n14657), .Y(n14649) );
  AOI21X1 U13824 ( .A(n14617), .B(\regX[21][6] ), .C(n14658), .Y(n14657) );
  OAI22X1 U13825 ( .A(n12849), .B(n14619), .C(n13173), .D(n14620), .Y(n14658)
         );
  INVX1 U13826 ( .A(\regX[23][6] ), .Y(n12849) );
  AOI22X1 U13827 ( .A(n14621), .B(N1683), .C(n14622), .D(\regX[19][6] ), .Y(
        n14656) );
  AOI22X1 U13828 ( .A(n14623), .B(\regX[13][6] ), .C(n14624), .D(\regX[20][6] ), .Y(n14655) );
  NOR2X1 U13829 ( .A(n14659), .B(n14660), .Y(n14647) );
  OAI21X1 U13830 ( .A(n12602), .B(n14627), .C(n14661), .Y(n14660) );
  AOI22X1 U13831 ( .A(n14629), .B(\regX[22][6] ), .C(n14630), .D(\regX[1][6] ), 
        .Y(n14661) );
  INVX1 U13832 ( .A(\regX[0][6] ), .Y(n12602) );
  OR2X1 U13833 ( .A(n14662), .B(n14663), .Y(n14659) );
  OAI22X1 U13834 ( .A(n12767), .B(n14633), .C(n12778), .D(n14634), .Y(n14663)
         );
  OAI21X1 U13835 ( .A(n12754), .B(n14635), .C(n12506), .Y(n14662) );
  NAND2X1 U13836 ( .A(N2752), .B(n15377), .Y(n12506) );
  INVX1 U13837 ( .A(\regX[7][6] ), .Y(n12754) );
  NOR2X1 U13838 ( .A(n14664), .B(n14665), .Y(n14646) );
  OAI21X1 U13839 ( .A(n12719), .B(n14638), .C(n14666), .Y(n14665) );
  AOI22X1 U13840 ( .A(n14640), .B(N1381), .C(\regX[6][6] ), .D(n14641), .Y(
        n14666) );
  OAI21X1 U13841 ( .A(n12898), .B(n14642), .C(n14667), .Y(n14664) );
  AOI22X1 U13842 ( .A(n14644), .B(\regX[5][6] ), .C(n14645), .D(N1621), .Y(
        n14667) );
  INVX1 U13843 ( .A(\regX[11][6] ), .Y(n12898) );
  NAND3X1 U13844 ( .A(n14668), .B(n14669), .C(n14670), .Y(\U3/U119/Z_5 ) );
  NOR2X1 U13845 ( .A(n14671), .B(n14672), .Y(n14670) );
  OR2X1 U13846 ( .A(n14673), .B(n14674), .Y(n14672) );
  OAI21X1 U13847 ( .A(n12799), .B(n14606), .C(n14675), .Y(n14674) );
  AOI22X1 U13848 ( .A(n14608), .B(\regX[16][5] ), .C(n14609), .D(\regX[24][5] ), .Y(n14675) );
  INVX1 U13849 ( .A(\regX[17][5] ), .Y(n12799) );
  OAI21X1 U13850 ( .A(n12730), .B(n14610), .C(n14676), .Y(n14673) );
  AOI22X1 U13851 ( .A(n14612), .B(\regX[15][5] ), .C(n14613), .D(N1740), .Y(
        n14676) );
  INVX1 U13852 ( .A(N1438), .Y(n12730) );
  NAND3X1 U13853 ( .A(n14677), .B(n14678), .C(n14679), .Y(n14671) );
  AOI21X1 U13854 ( .A(n14617), .B(\regX[21][5] ), .C(n14680), .Y(n14679) );
  OAI22X1 U13855 ( .A(n12848), .B(n14619), .C(n13172), .D(n14620), .Y(n14680)
         );
  INVX1 U13856 ( .A(\regX[23][5] ), .Y(n12848) );
  AOI22X1 U13857 ( .A(n14621), .B(N1682), .C(n14622), .D(\regX[19][5] ), .Y(
        n14678) );
  AOI22X1 U13858 ( .A(n14623), .B(\regX[13][5] ), .C(n14624), .D(\regX[20][5] ), .Y(n14677) );
  NOR2X1 U13859 ( .A(n14681), .B(n14682), .Y(n14669) );
  OAI21X1 U13860 ( .A(n12601), .B(n14627), .C(n14683), .Y(n14682) );
  AOI22X1 U13861 ( .A(n14629), .B(\regX[22][5] ), .C(n14630), .D(\regX[1][5] ), 
        .Y(n14683) );
  INVX1 U13862 ( .A(\regX[0][5] ), .Y(n12601) );
  OR2X1 U13863 ( .A(n14684), .B(n14685), .Y(n14681) );
  OAI22X1 U13864 ( .A(n12766), .B(n14633), .C(n12777), .D(n14634), .Y(n14685)
         );
  OAI21X1 U13865 ( .A(n12753), .B(n14635), .C(n12507), .Y(n14684) );
  NAND2X1 U13866 ( .A(N2751), .B(n15377), .Y(n12507) );
  INVX1 U13867 ( .A(\regX[7][5] ), .Y(n12753) );
  NOR2X1 U13868 ( .A(n14686), .B(n14687), .Y(n14668) );
  OAI21X1 U13869 ( .A(n12718), .B(n14638), .C(n14688), .Y(n14687) );
  AOI22X1 U13870 ( .A(n14640), .B(N1380), .C(\regX[6][5] ), .D(n14641), .Y(
        n14688) );
  OAI21X1 U13871 ( .A(n12897), .B(n14642), .C(n14689), .Y(n14686) );
  AOI22X1 U13872 ( .A(n14644), .B(\regX[5][5] ), .C(n14645), .D(N1620), .Y(
        n14689) );
  INVX1 U13873 ( .A(\regX[11][5] ), .Y(n12897) );
  NAND3X1 U13874 ( .A(n14690), .B(n14691), .C(n14692), .Y(\U3/U119/Z_4 ) );
  NOR2X1 U13875 ( .A(n14693), .B(n14694), .Y(n14692) );
  OR2X1 U13876 ( .A(n14695), .B(n14696), .Y(n14694) );
  OAI21X1 U13877 ( .A(n12798), .B(n14606), .C(n14697), .Y(n14696) );
  AOI22X1 U13878 ( .A(n14608), .B(\regX[16][4] ), .C(n14609), .D(\regX[24][4] ), .Y(n14697) );
  INVX1 U13879 ( .A(n14698), .Y(n14608) );
  INVX1 U13880 ( .A(\regX[17][4] ), .Y(n12798) );
  OAI21X1 U13881 ( .A(n12729), .B(n14610), .C(n14699), .Y(n14695) );
  AOI22X1 U13882 ( .A(n14612), .B(\regX[15][4] ), .C(n14613), .D(N1739), .Y(
        n14699) );
  INVX1 U13883 ( .A(N1437), .Y(n12729) );
  NAND3X1 U13884 ( .A(n14700), .B(n14701), .C(n14702), .Y(n14693) );
  AOI21X1 U13885 ( .A(n14617), .B(\regX[21][4] ), .C(n14703), .Y(n14702) );
  OAI22X1 U13886 ( .A(n12847), .B(n14619), .C(n13171), .D(n14620), .Y(n14703)
         );
  INVX1 U13887 ( .A(\regX[23][4] ), .Y(n12847) );
  INVX1 U13888 ( .A(n14704), .Y(n14617) );
  AOI22X1 U13889 ( .A(n14621), .B(N1681), .C(n14622), .D(\regX[19][4] ), .Y(
        n14701) );
  INVX1 U13890 ( .A(n14705), .Y(n14621) );
  AOI22X1 U13891 ( .A(n14623), .B(\regX[13][4] ), .C(n14624), .D(\regX[20][4] ), .Y(n14700) );
  NOR2X1 U13892 ( .A(n14706), .B(n14707), .Y(n14691) );
  OAI21X1 U13893 ( .A(n12600), .B(n14627), .C(n14708), .Y(n14707) );
  AOI22X1 U13894 ( .A(n14629), .B(\regX[22][4] ), .C(n14630), .D(\regX[1][4] ), 
        .Y(n14708) );
  INVX1 U13895 ( .A(\regX[0][4] ), .Y(n12600) );
  OR2X1 U13896 ( .A(n14709), .B(n14710), .Y(n14706) );
  OAI22X1 U13897 ( .A(n12765), .B(n14633), .C(n12776), .D(n14634), .Y(n14710)
         );
  OAI21X1 U13898 ( .A(n12752), .B(n14635), .C(n12508), .Y(n14709) );
  NAND2X1 U13899 ( .A(N2750), .B(n15377), .Y(n12508) );
  INVX1 U13900 ( .A(\regX[7][4] ), .Y(n12752) );
  NOR2X1 U13901 ( .A(n14711), .B(n14712), .Y(n14690) );
  OAI21X1 U13902 ( .A(n12717), .B(n14638), .C(n14713), .Y(n14712) );
  AOI22X1 U13903 ( .A(n14640), .B(N1379), .C(\regX[6][4] ), .D(n14641), .Y(
        n14713) );
  INVX1 U13904 ( .A(n14714), .Y(n14640) );
  OAI21X1 U13905 ( .A(n12896), .B(n14642), .C(n14715), .Y(n14711) );
  AOI22X1 U13906 ( .A(n14644), .B(\regX[5][4] ), .C(n14645), .D(N1619), .Y(
        n14715) );
  INVX1 U13907 ( .A(n14716), .Y(n14644) );
  INVX1 U13908 ( .A(\regX[11][4] ), .Y(n12896) );
  NOR2X1 U13909 ( .A(n14214), .B(n13032), .Y(\U3/U119/Z_31 ) );
  INVX1 U13910 ( .A(N2776), .Y(n13032) );
  NAND3X1 U13911 ( .A(n14717), .B(n14718), .C(n14719), .Y(\U3/U119/Z_3 ) );
  NOR2X1 U13912 ( .A(n14720), .B(n14721), .Y(n14719) );
  OR2X1 U13913 ( .A(n14722), .B(n14723), .Y(n14721) );
  OAI21X1 U13914 ( .A(n14214), .B(n14295), .C(n14724), .Y(n14723) );
  AOI22X1 U13915 ( .A(n14609), .B(\regX[24][3] ), .C(n14725), .D(\regX[17][3] ), .Y(n14724) );
  OAI21X1 U13916 ( .A(n12786), .B(n14698), .C(n14726), .Y(n14722) );
  AOI22X1 U13917 ( .A(n14613), .B(N1738), .C(n14727), .D(N1436), .Y(n14726) );
  INVX1 U13918 ( .A(\regX[16][3] ), .Y(n12786) );
  NAND3X1 U13919 ( .A(n14728), .B(n14729), .C(n14730), .Y(n14720) );
  AOI21X1 U13920 ( .A(n14612), .B(\regX[15][3] ), .C(n14731), .Y(n14730) );
  OAI22X1 U13921 ( .A(n12875), .B(n14704), .C(n12846), .D(n14619), .Y(n14731)
         );
  INVX1 U13922 ( .A(\regX[23][3] ), .Y(n12846) );
  AOI22X1 U13923 ( .A(n14622), .B(\regX[19][3] ), .C(n14623), .D(\regX[13][3] ), .Y(n14729) );
  AOI22X1 U13924 ( .A(n14624), .B(\regX[20][3] ), .C(n14732), .D(\regX[18][3] ), .Y(n14728) );
  NOR2X1 U13925 ( .A(n14733), .B(n14734), .Y(n14718) );
  OAI21X1 U13926 ( .A(n12740), .B(n14716), .C(n14735), .Y(n14734) );
  AOI22X1 U13927 ( .A(n14630), .B(\regX[1][3] ), .C(n14736), .D(\regX[0][3] ), 
        .Y(n14735) );
  INVX1 U13928 ( .A(\regX[5][3] ), .Y(n12740) );
  NAND2X1 U13929 ( .A(n14737), .B(n14738), .Y(n14733) );
  AOI22X1 U13930 ( .A(n14739), .B(\regX[7][3] ), .C(n14740), .D(\regX[9][3] ), 
        .Y(n14738) );
  AOI22X1 U13931 ( .A(n14741), .B(\regX[8][3] ), .C(n14629), .D(\regX[22][3] ), 
        .Y(n14737) );
  NOR2X1 U13932 ( .A(n14742), .B(n14743), .Y(n14717) );
  OAI21X1 U13933 ( .A(n12856), .B(n14705), .C(n14744), .Y(n14743) );
  AOI22X1 U13934 ( .A(\regX[6][3] ), .B(n14641), .C(n14745), .D(\regX[3][3] ), 
        .Y(n14744) );
  OAI21X1 U13935 ( .A(n12705), .B(n14714), .C(n14746), .Y(n14742) );
  AOI22X1 U13936 ( .A(n14645), .B(N1618), .C(n14747), .D(\regX[11][3] ), .Y(
        n14746) );
  NOR2X1 U13937 ( .A(n14214), .B(n14296), .Y(\U3/U119/Z_29 ) );
  INVX1 U13938 ( .A(N2775), .Y(n14296) );
  NOR2X1 U13939 ( .A(n14214), .B(n14298), .Y(\U3/U119/Z_28 ) );
  INVX1 U13940 ( .A(N2774), .Y(n14298) );
  NOR2X1 U13941 ( .A(n14214), .B(n14299), .Y(\U3/U119/Z_27 ) );
  INVX1 U13942 ( .A(N2773), .Y(n14299) );
  NOR2X1 U13943 ( .A(n14214), .B(n14300), .Y(\U3/U119/Z_26 ) );
  INVX1 U13944 ( .A(N2772), .Y(n14300) );
  NOR2X1 U13945 ( .A(n14214), .B(n14301), .Y(\U3/U119/Z_25 ) );
  INVX1 U13946 ( .A(N2771), .Y(n14301) );
  NOR2X1 U13947 ( .A(n14214), .B(n14302), .Y(\U3/U119/Z_24 ) );
  INVX1 U13948 ( .A(N2770), .Y(n14302) );
  NOR2X1 U13949 ( .A(n14214), .B(n14303), .Y(\U3/U119/Z_23 ) );
  INVX1 U13950 ( .A(N2769), .Y(n14303) );
  NOR2X1 U13951 ( .A(n14214), .B(n14304), .Y(\U3/U119/Z_22 ) );
  INVX1 U13952 ( .A(N2768), .Y(n14304) );
  NOR2X1 U13953 ( .A(n14214), .B(n14305), .Y(\U3/U119/Z_21 ) );
  INVX1 U13954 ( .A(N2767), .Y(n14305) );
  NOR2X1 U13955 ( .A(n14214), .B(n14306), .Y(\U3/U119/Z_20 ) );
  INVX1 U13956 ( .A(N2766), .Y(n14306) );
  NAND3X1 U13957 ( .A(n14748), .B(n14749), .C(n14750), .Y(\U3/U119/Z_2 ) );
  NOR2X1 U13958 ( .A(n14751), .B(n14752), .Y(n14750) );
  OR2X1 U13959 ( .A(n14753), .B(n14754), .Y(n14752) );
  OAI21X1 U13960 ( .A(n14214), .B(n14297), .C(n14755), .Y(n14754) );
  AOI22X1 U13961 ( .A(n14609), .B(\regX[24][2] ), .C(n14725), .D(\regX[17][2] ), .Y(n14755) );
  OAI21X1 U13962 ( .A(n12785), .B(n14698), .C(n14756), .Y(n14753) );
  AOI22X1 U13963 ( .A(n14613), .B(N1737), .C(n14727), .D(N1435), .Y(n14756) );
  INVX1 U13964 ( .A(\regX[16][2] ), .Y(n12785) );
  NAND3X1 U13965 ( .A(n14757), .B(n14758), .C(n14759), .Y(n14751) );
  AOI21X1 U13966 ( .A(n14612), .B(\regX[15][2] ), .C(n14760), .Y(n14759) );
  OAI22X1 U13967 ( .A(n12874), .B(n14704), .C(n12845), .D(n14619), .Y(n14760)
         );
  INVX1 U13968 ( .A(\regX[23][2] ), .Y(n12845) );
  AOI22X1 U13969 ( .A(n14622), .B(\regX[19][2] ), .C(n14623), .D(\regX[13][2] ), .Y(n14758) );
  AOI22X1 U13970 ( .A(n14624), .B(\regX[20][2] ), .C(n14732), .D(\regX[18][2] ), .Y(n14757) );
  NOR2X1 U13971 ( .A(n14761), .B(n14762), .Y(n14749) );
  OAI21X1 U13972 ( .A(n12739), .B(n14716), .C(n14763), .Y(n14762) );
  AOI22X1 U13973 ( .A(n14630), .B(\regX[1][2] ), .C(n14736), .D(\regX[0][2] ), 
        .Y(n14763) );
  INVX1 U13974 ( .A(\regX[5][2] ), .Y(n12739) );
  NAND2X1 U13975 ( .A(n14764), .B(n14765), .Y(n14761) );
  AOI22X1 U13976 ( .A(n14739), .B(\regX[7][2] ), .C(n14740), .D(\regX[9][2] ), 
        .Y(n14765) );
  AOI22X1 U13977 ( .A(n14741), .B(\regX[8][2] ), .C(n14629), .D(\regX[22][2] ), 
        .Y(n14764) );
  NOR2X1 U13978 ( .A(n14766), .B(n14767), .Y(n14748) );
  OAI21X1 U13979 ( .A(n12855), .B(n14705), .C(n14768), .Y(n14767) );
  AOI22X1 U13980 ( .A(\regX[6][2] ), .B(n14641), .C(n14745), .D(\regX[3][2] ), 
        .Y(n14768) );
  OAI21X1 U13981 ( .A(n12704), .B(n14714), .C(n14769), .Y(n14766) );
  AOI22X1 U13982 ( .A(n14645), .B(N1617), .C(n14747), .D(\regX[11][2] ), .Y(
        n14769) );
  NOR2X1 U13983 ( .A(n14214), .B(n14307), .Y(\U3/U119/Z_19 ) );
  INVX1 U13984 ( .A(N2765), .Y(n14307) );
  NOR2X1 U13985 ( .A(n14214), .B(n14309), .Y(\U3/U119/Z_18 ) );
  INVX1 U13986 ( .A(N2764), .Y(n14309) );
  NOR2X1 U13987 ( .A(n14214), .B(n14310), .Y(\U3/U119/Z_17 ) );
  INVX1 U13988 ( .A(N2763), .Y(n14310) );
  NOR2X1 U13989 ( .A(n14214), .B(n14311), .Y(\U3/U119/Z_16 ) );
  INVX1 U13990 ( .A(N2762), .Y(n14311) );
  NOR2X1 U13991 ( .A(n14214), .B(n14312), .Y(\U3/U119/Z_15 ) );
  INVX1 U13992 ( .A(N2761), .Y(n14312) );
  NOR2X1 U13993 ( .A(n14214), .B(n14313), .Y(\U3/U119/Z_14 ) );
  INVX1 U13994 ( .A(N2760), .Y(n14313) );
  NOR2X1 U13995 ( .A(n14214), .B(n14314), .Y(\U3/U119/Z_13 ) );
  INVX1 U13996 ( .A(N2759), .Y(n14314) );
  NOR2X1 U13997 ( .A(n14214), .B(n14315), .Y(\U3/U119/Z_12 ) );
  INVX1 U13998 ( .A(N2758), .Y(n14315) );
  NOR2X1 U13999 ( .A(n14214), .B(n14316), .Y(\U3/U119/Z_11 ) );
  INVX1 U14000 ( .A(N2757), .Y(n14316) );
  NOR2X1 U14001 ( .A(n14214), .B(n14317), .Y(\U3/U119/Z_10 ) );
  INVX1 U14002 ( .A(N2756), .Y(n14317) );
  NAND3X1 U14003 ( .A(n14770), .B(n14771), .C(n14772), .Y(\U3/U119/Z_1 ) );
  NOR2X1 U14004 ( .A(n14773), .B(n14774), .Y(n14772) );
  OR2X1 U14005 ( .A(n14775), .B(n14776), .Y(n14774) );
  OAI21X1 U14006 ( .A(n14214), .B(n14308), .C(n14777), .Y(n14776) );
  AOI22X1 U14007 ( .A(n14609), .B(\regX[24][1] ), .C(n14725), .D(\regX[17][1] ), .Y(n14777) );
  OAI21X1 U14008 ( .A(n12784), .B(n14698), .C(n14778), .Y(n14775) );
  AOI22X1 U14009 ( .A(n14613), .B(N1736), .C(n14727), .D(N1434), .Y(n14778) );
  INVX1 U14010 ( .A(\regX[16][1] ), .Y(n12784) );
  NAND3X1 U14011 ( .A(n14779), .B(n14780), .C(n14781), .Y(n14773) );
  AOI21X1 U14012 ( .A(n14612), .B(\regX[15][1] ), .C(n14782), .Y(n14781) );
  OAI22X1 U14013 ( .A(n12873), .B(n14704), .C(n12844), .D(n14619), .Y(n14782)
         );
  INVX1 U14014 ( .A(\regX[23][1] ), .Y(n12844) );
  AOI22X1 U14015 ( .A(n14622), .B(\regX[19][1] ), .C(n14623), .D(\regX[13][1] ), .Y(n14780) );
  AOI22X1 U14016 ( .A(n14624), .B(\regX[20][1] ), .C(n14732), .D(\regX[18][1] ), .Y(n14779) );
  NOR2X1 U14017 ( .A(n14783), .B(n14784), .Y(n14771) );
  OAI21X1 U14018 ( .A(n12738), .B(n14716), .C(n14785), .Y(n14784) );
  AOI22X1 U14019 ( .A(n14630), .B(\regX[1][1] ), .C(n14736), .D(\regX[0][1] ), 
        .Y(n14785) );
  INVX1 U14020 ( .A(\regX[5][1] ), .Y(n12738) );
  NAND2X1 U14021 ( .A(n14786), .B(n14787), .Y(n14783) );
  AOI22X1 U14022 ( .A(n14739), .B(\regX[7][1] ), .C(n14740), .D(\regX[9][1] ), 
        .Y(n14787) );
  AOI22X1 U14023 ( .A(n14741), .B(\regX[8][1] ), .C(n14629), .D(\regX[22][1] ), 
        .Y(n14786) );
  NOR2X1 U14024 ( .A(n14788), .B(n14789), .Y(n14770) );
  OAI21X1 U14025 ( .A(n12854), .B(n14705), .C(n14790), .Y(n14789) );
  AOI22X1 U14026 ( .A(\regX[6][1] ), .B(n14641), .C(n14745), .D(\regX[3][1] ), 
        .Y(n14790) );
  OAI21X1 U14027 ( .A(n12703), .B(n14714), .C(n14791), .Y(n14788) );
  AOI22X1 U14028 ( .A(n14645), .B(N1616), .C(n14747), .D(\regX[11][1] ), .Y(
        n14791) );
  NAND3X1 U14029 ( .A(n14792), .B(n14793), .C(n14794), .Y(\U3/U119/Z_0 ) );
  NOR2X1 U14030 ( .A(n14795), .B(n14796), .Y(n14794) );
  OR2X1 U14031 ( .A(n14797), .B(n14798), .Y(n14796) );
  OAI21X1 U14032 ( .A(n14214), .B(n14319), .C(n14799), .Y(n14798) );
  AOI22X1 U14033 ( .A(n14609), .B(\regX[24][0] ), .C(n14725), .D(\regX[17][0] ), .Y(n14799) );
  INVX1 U14034 ( .A(n14606), .Y(n14725) );
  NAND2X1 U14035 ( .A(n14800), .B(n14801), .Y(n14606) );
  AND2X1 U14036 ( .A(n14802), .B(n14803), .Y(n14609) );
  OAI21X1 U14037 ( .A(n12782), .B(n14698), .C(n14804), .Y(n14797) );
  AOI22X1 U14038 ( .A(n14613), .B(N1735), .C(n14727), .D(N1433), .Y(n14804) );
  INVX1 U14039 ( .A(n14610), .Y(n14727) );
  NAND2X1 U14040 ( .A(n14805), .B(n14806), .Y(n14610) );
  AND2X1 U14041 ( .A(n14807), .B(n14808), .Y(n14613) );
  NAND3X1 U14042 ( .A(n14809), .B(n14801), .C(n14810), .Y(n14698) );
  INVX1 U14043 ( .A(\regX[16][0] ), .Y(n12782) );
  NAND3X1 U14044 ( .A(n14811), .B(n14812), .C(n14813), .Y(n14795) );
  AOI21X1 U14045 ( .A(n14612), .B(\regX[15][0] ), .C(n14814), .Y(n14813) );
  OAI22X1 U14046 ( .A(n12871), .B(n14704), .C(n12842), .D(n14619), .Y(n14814)
         );
  NAND2X1 U14047 ( .A(n14800), .B(n14808), .Y(n14619) );
  INVX1 U14048 ( .A(\regX[23][0] ), .Y(n12842) );
  NAND2X1 U14049 ( .A(n14800), .B(n14805), .Y(n14704) );
  AND2X1 U14050 ( .A(n14815), .B(n14808), .Y(n14612) );
  AOI22X1 U14051 ( .A(n14622), .B(\regX[19][0] ), .C(n14623), .D(\regX[13][0] ), .Y(n14812) );
  AND2X1 U14052 ( .A(n14805), .B(n14815), .Y(n14623) );
  AND2X1 U14053 ( .A(n14800), .B(n14816), .Y(n14622) );
  INVX1 U14054 ( .A(n14817), .Y(n14800) );
  NAND3X1 U14055 ( .A(n15328), .B(n14803), .C(n14818), .Y(n14817) );
  AOI22X1 U14056 ( .A(n14624), .B(\regX[20][0] ), .C(n14732), .D(\regX[18][0] ), .Y(n14811) );
  INVX1 U14057 ( .A(n14620), .Y(n14732) );
  NAND2X1 U14058 ( .A(n14816), .B(n14810), .Y(n14620) );
  AND2X1 U14059 ( .A(n14805), .B(n14810), .Y(n14624) );
  NOR2X1 U14060 ( .A(n14819), .B(n14820), .Y(n14793) );
  OAI21X1 U14061 ( .A(n12736), .B(n14716), .C(n14821), .Y(n14820) );
  AOI22X1 U14062 ( .A(n14630), .B(\regX[1][0] ), .C(n14736), .D(\regX[0][0] ), 
        .Y(n14821) );
  INVX1 U14063 ( .A(n14627), .Y(n14736) );
  NAND2X1 U14064 ( .A(n14806), .B(n14801), .Y(n14627) );
  AND2X1 U14065 ( .A(n14801), .B(n14822), .Y(n14630) );
  NAND2X1 U14066 ( .A(n14805), .B(n14822), .Y(n14716) );
  INVX1 U14067 ( .A(\regX[5][0] ), .Y(n12736) );
  NAND2X1 U14068 ( .A(n14823), .B(n14824), .Y(n14819) );
  AOI22X1 U14069 ( .A(n14739), .B(\regX[7][0] ), .C(n14740), .D(\regX[9][0] ), 
        .Y(n14824) );
  INVX1 U14070 ( .A(n14634), .Y(n14740) );
  NAND2X1 U14071 ( .A(n14801), .B(n14815), .Y(n14634) );
  INVX1 U14072 ( .A(n14635), .Y(n14739) );
  NAND2X1 U14073 ( .A(n14808), .B(n14822), .Y(n14635) );
  AOI22X1 U14074 ( .A(n14741), .B(\regX[8][0] ), .C(n14629), .D(\regX[22][0] ), 
        .Y(n14823) );
  AND2X1 U14075 ( .A(n14810), .B(n14808), .Y(n14629) );
  INVX1 U14076 ( .A(n14825), .Y(n14810) );
  NAND3X1 U14077 ( .A(n14803), .B(n14826), .C(n15328), .Y(n14825) );
  INVX1 U14078 ( .A(n14633), .Y(n14741) );
  NAND3X1 U14079 ( .A(n14827), .B(n14801), .C(n14807), .Y(n14633) );
  NOR2X1 U14080 ( .A(n14828), .B(n14829), .Y(n14801) );
  NOR2X1 U14081 ( .A(n14830), .B(n14831), .Y(n14792) );
  OAI21X1 U14082 ( .A(n12852), .B(n14705), .C(n14832), .Y(n14831) );
  AOI22X1 U14083 ( .A(\regX[6][0] ), .B(n14641), .C(n14745), .D(\regX[3][0] ), 
        .Y(n14832) );
  INVX1 U14084 ( .A(n14638), .Y(n14745) );
  NAND2X1 U14085 ( .A(n14816), .B(n14822), .Y(n14638) );
  NOR2X1 U14086 ( .A(n14833), .B(n14826), .Y(n14822) );
  INVX1 U14087 ( .A(n14834), .Y(n14641) );
  AOI21X1 U14088 ( .A(n14808), .B(n14806), .C(n15369), .Y(n14834) );
  NOR2X1 U14089 ( .A(n14835), .B(n14836), .Y(n14808) );
  NAND2X1 U14090 ( .A(n14805), .B(n14807), .Y(n14705) );
  NOR2X1 U14091 ( .A(n14829), .B(n14835), .Y(n14805) );
  INVX1 U14092 ( .A(n14828), .Y(n14835) );
  OAI21X1 U14093 ( .A(n12701), .B(n14714), .C(n14837), .Y(n14830) );
  AOI22X1 U14094 ( .A(n14645), .B(N1615), .C(n14747), .D(\regX[11][0] ), .Y(
        n14837) );
  INVX1 U14095 ( .A(n14642), .Y(n14747) );
  NAND2X1 U14096 ( .A(n14816), .B(n14815), .Y(n14642) );
  AND2X1 U14097 ( .A(n14802), .B(n14818), .Y(n14815) );
  AND2X1 U14098 ( .A(n14816), .B(n14807), .Y(n14645) );
  AND2X1 U14099 ( .A(n14802), .B(n14826), .Y(n14807) );
  NOR2X1 U14100 ( .A(n14809), .B(n12552), .Y(n14802) );
  NAND2X1 U14101 ( .A(n14816), .B(n14806), .Y(n14714) );
  NOR2X1 U14102 ( .A(n14833), .B(n14818), .Y(n14806) );
  NAND3X1 U14103 ( .A(n14809), .B(n15328), .C(n14827), .Y(n14833) );
  INVX1 U14104 ( .A(n14803), .Y(n14827) );
  XOR2X1 U14105 ( .A(n14838), .B(n14839), .Y(n14803) );
  XOR2X1 U14106 ( .A(n14840), .B(n14841), .Y(n14839) );
  OAI21X1 U14107 ( .A(n14842), .B(n14843), .C(n14844), .Y(n14841) );
  OAI21X1 U14108 ( .A(n14845), .B(n14846), .C(n14582), .Y(n14844) );
  AND2X1 U14109 ( .A(N3343), .B(n15328), .Y(n14582) );
  OR2X1 U14110 ( .A(n14845), .B(N3343), .Y(n14843) );
  INVX1 U14111 ( .A(n14847), .Y(n14842) );
  OAI21X1 U14112 ( .A(n14848), .B(n14849), .C(n14850), .Y(n14840) );
  OAI21X1 U14113 ( .A(n14851), .B(n14852), .C(n14838), .Y(n14850) );
  INVX1 U14114 ( .A(n14849), .Y(n14852) );
  NOR2X1 U14115 ( .A(n14828), .B(n14836), .Y(n14816) );
  INVX1 U14116 ( .A(n14829), .Y(n14836) );
  NOR2X1 U14117 ( .A(n14214), .B(n12986), .Y(\U3/U118/Z_9 ) );
  INVX1 U14118 ( .A(fGy[9]), .Y(n12986) );
  NOR2X1 U14119 ( .A(n14214), .B(n12984), .Y(\U3/U118/Z_8 ) );
  INVX1 U14120 ( .A(fGy[8]), .Y(n12984) );
  OAI21X1 U14121 ( .A(n14853), .B(n13921), .C(n12514), .Y(\U3/U118/Z_7 ) );
  NAND2X1 U14122 ( .A(fGy[7]), .B(n15377), .Y(n12514) );
  NOR2X1 U14123 ( .A(n14854), .B(n14855), .Y(n14853) );
  NAND2X1 U14124 ( .A(n14856), .B(n14857), .Y(n14855) );
  NOR2X1 U14125 ( .A(n14858), .B(n14859), .Y(n14857) );
  OAI21X1 U14126 ( .A(n12677), .B(n14860), .C(n14861), .Y(n14859) );
  AOI22X1 U14127 ( .A(n14862), .B(\regX[11][7] ), .C(n14863), .D(\regX[7][7] ), 
        .Y(n14861) );
  OAI21X1 U14128 ( .A(n12698), .B(n14864), .C(n14865), .Y(n14858) );
  AOI22X1 U14129 ( .A(n14866), .B(N1622), .C(n14867), .D(\regX[23][7] ), .Y(
        n14865) );
  INVX1 U14130 ( .A(\regX[1][7] ), .Y(n12698) );
  NOR2X1 U14131 ( .A(n14868), .B(n14869), .Y(n14856) );
  OAI21X1 U14132 ( .A(n12779), .B(n14870), .C(n14871), .Y(n14869) );
  AOI22X1 U14133 ( .A(n14872), .B(\regX[5][7] ), .C(n14873), .D(\regX[0][7] ), 
        .Y(n14871) );
  INVX1 U14134 ( .A(\regX[9][7] ), .Y(n12779) );
  OAI21X1 U14135 ( .A(n12709), .B(n14874), .C(n14875), .Y(n14868) );
  AOI22X1 U14136 ( .A(n14876), .B(\regX[13][7] ), .C(n14877), .D(N1440), .Y(
        n14875) );
  NAND3X1 U14137 ( .A(n14878), .B(n14879), .C(n14880), .Y(n14854) );
  NOR2X1 U14138 ( .A(n14881), .B(n14882), .Y(n14880) );
  OAI21X1 U14139 ( .A(n12768), .B(n14883), .C(n14884), .Y(n14882) );
  AOI22X1 U14140 ( .A(n14885), .B(N1684), .C(n14886), .D(\regX[17][7] ), .Y(
        n14884) );
  INVX1 U14141 ( .A(\regX[8][7] ), .Y(n12768) );
  OAI21X1 U14142 ( .A(n12591), .B(n14887), .C(n14888), .Y(n14881) );
  AOI22X1 U14143 ( .A(n14889), .B(N1742), .C(n14890), .D(\regX[19][7] ), .Y(
        n14888) );
  INVX1 U14144 ( .A(\regX[15][7] ), .Y(n12591) );
  NOR2X1 U14145 ( .A(n14891), .B(n14892), .Y(n14879) );
  OAI22X1 U14146 ( .A(n12720), .B(n14893), .C(n12840), .D(n14894), .Y(n14892)
         );
  INVX1 U14147 ( .A(\regX[22][7] ), .Y(n12840) );
  INVX1 U14148 ( .A(\regX[3][7] ), .Y(n12720) );
  OAI22X1 U14149 ( .A(n12869), .B(n14895), .C(n12812), .D(n14896), .Y(n14891)
         );
  INVX1 U14150 ( .A(\regX[24][7] ), .Y(n12812) );
  INVX1 U14151 ( .A(\regX[20][7] ), .Y(n12869) );
  AOI21X1 U14152 ( .A(n14897), .B(\regX[16][7] ), .C(n14898), .Y(n14878) );
  OAI22X1 U14153 ( .A(n13174), .B(n14899), .C(n12879), .D(n14900), .Y(n14898)
         );
  INVX1 U14154 ( .A(\regX[21][7] ), .Y(n12879) );
  OAI21X1 U14155 ( .A(n14901), .B(n13921), .C(n12515), .Y(\U3/U118/Z_6 ) );
  NAND2X1 U14156 ( .A(fGy[6]), .B(n15377), .Y(n12515) );
  NOR2X1 U14157 ( .A(n14902), .B(n14903), .Y(n14901) );
  NAND2X1 U14158 ( .A(n14904), .B(n14905), .Y(n14903) );
  NOR2X1 U14159 ( .A(n14906), .B(n14907), .Y(n14905) );
  OAI21X1 U14160 ( .A(n12676), .B(n14860), .C(n14908), .Y(n14907) );
  AOI22X1 U14161 ( .A(n14862), .B(\regX[11][6] ), .C(n14863), .D(\regX[7][6] ), 
        .Y(n14908) );
  OAI21X1 U14162 ( .A(n12697), .B(n14864), .C(n14909), .Y(n14906) );
  AOI22X1 U14163 ( .A(n14866), .B(N1621), .C(n14867), .D(\regX[23][6] ), .Y(
        n14909) );
  INVX1 U14164 ( .A(\regX[1][6] ), .Y(n12697) );
  NOR2X1 U14165 ( .A(n14910), .B(n14911), .Y(n14904) );
  OAI21X1 U14166 ( .A(n12778), .B(n14870), .C(n14912), .Y(n14911) );
  AOI22X1 U14167 ( .A(n14872), .B(\regX[5][6] ), .C(n14873), .D(\regX[0][6] ), 
        .Y(n14912) );
  INVX1 U14168 ( .A(\regX[9][6] ), .Y(n12778) );
  OAI21X1 U14169 ( .A(n12708), .B(n14874), .C(n14913), .Y(n14910) );
  AOI22X1 U14170 ( .A(n14876), .B(\regX[13][6] ), .C(n14877), .D(N1439), .Y(
        n14913) );
  NAND3X1 U14171 ( .A(n14914), .B(n14915), .C(n14916), .Y(n14902) );
  NOR2X1 U14172 ( .A(n14917), .B(n14918), .Y(n14916) );
  OAI21X1 U14173 ( .A(n12767), .B(n14883), .C(n14919), .Y(n14918) );
  AOI22X1 U14174 ( .A(n14885), .B(N1683), .C(n14886), .D(\regX[17][6] ), .Y(
        n14919) );
  INVX1 U14175 ( .A(\regX[8][6] ), .Y(n12767) );
  OAI21X1 U14176 ( .A(n12589), .B(n14887), .C(n14920), .Y(n14917) );
  AOI22X1 U14177 ( .A(n14889), .B(N1741), .C(n14890), .D(\regX[19][6] ), .Y(
        n14920) );
  INVX1 U14178 ( .A(\regX[15][6] ), .Y(n12589) );
  NOR2X1 U14179 ( .A(n14921), .B(n14922), .Y(n14915) );
  OAI22X1 U14180 ( .A(n12719), .B(n14893), .C(n12839), .D(n14894), .Y(n14922)
         );
  INVX1 U14181 ( .A(\regX[22][6] ), .Y(n12839) );
  INVX1 U14182 ( .A(\regX[3][6] ), .Y(n12719) );
  OAI22X1 U14183 ( .A(n12868), .B(n14895), .C(n12811), .D(n14896), .Y(n14921)
         );
  INVX1 U14184 ( .A(\regX[24][6] ), .Y(n12811) );
  INVX1 U14185 ( .A(\regX[20][6] ), .Y(n12868) );
  AOI21X1 U14186 ( .A(n14897), .B(\regX[16][6] ), .C(n14923), .Y(n14914) );
  OAI22X1 U14187 ( .A(n13173), .B(n14899), .C(n12878), .D(n14900), .Y(n14923)
         );
  INVX1 U14188 ( .A(\regX[21][6] ), .Y(n12878) );
  OAI21X1 U14189 ( .A(n14924), .B(n13921), .C(n12516), .Y(\U3/U118/Z_5 ) );
  NAND2X1 U14190 ( .A(fGy[5]), .B(n15377), .Y(n12516) );
  NOR2X1 U14191 ( .A(n14925), .B(n14926), .Y(n14924) );
  NAND2X1 U14192 ( .A(n14927), .B(n14928), .Y(n14926) );
  NOR2X1 U14193 ( .A(n14929), .B(n14930), .Y(n14928) );
  OAI21X1 U14194 ( .A(n12675), .B(n14860), .C(n14931), .Y(n14930) );
  AOI22X1 U14195 ( .A(n14862), .B(\regX[11][5] ), .C(n14863), .D(\regX[7][5] ), 
        .Y(n14931) );
  INVX1 U14196 ( .A(\regX[6][5] ), .Y(n12675) );
  OAI21X1 U14197 ( .A(n12696), .B(n14864), .C(n14932), .Y(n14929) );
  AOI22X1 U14198 ( .A(n14866), .B(N1620), .C(n14867), .D(\regX[23][5] ), .Y(
        n14932) );
  INVX1 U14199 ( .A(\regX[1][5] ), .Y(n12696) );
  NOR2X1 U14200 ( .A(n14933), .B(n14934), .Y(n14927) );
  OAI21X1 U14201 ( .A(n12777), .B(n14870), .C(n14935), .Y(n14934) );
  AOI22X1 U14202 ( .A(n14872), .B(\regX[5][5] ), .C(n14873), .D(\regX[0][5] ), 
        .Y(n14935) );
  INVX1 U14203 ( .A(\regX[9][5] ), .Y(n12777) );
  OAI21X1 U14204 ( .A(n12707), .B(n14874), .C(n14936), .Y(n14933) );
  AOI22X1 U14205 ( .A(n14876), .B(\regX[13][5] ), .C(n14877), .D(N1438), .Y(
        n14936) );
  NAND3X1 U14206 ( .A(n14937), .B(n14938), .C(n14939), .Y(n14925) );
  NOR2X1 U14207 ( .A(n14940), .B(n14941), .Y(n14939) );
  OAI21X1 U14208 ( .A(n12766), .B(n14883), .C(n14942), .Y(n14941) );
  AOI22X1 U14209 ( .A(n14885), .B(N1682), .C(n14886), .D(\regX[17][5] ), .Y(
        n14942) );
  INVX1 U14210 ( .A(\regX[8][5] ), .Y(n12766) );
  OAI21X1 U14211 ( .A(n12587), .B(n14887), .C(n14943), .Y(n14940) );
  AOI22X1 U14212 ( .A(n14889), .B(N1740), .C(n14890), .D(\regX[19][5] ), .Y(
        n14943) );
  INVX1 U14213 ( .A(\regX[15][5] ), .Y(n12587) );
  NOR2X1 U14214 ( .A(n14944), .B(n14945), .Y(n14938) );
  OAI22X1 U14215 ( .A(n12718), .B(n14893), .C(n12838), .D(n14894), .Y(n14945)
         );
  INVX1 U14216 ( .A(\regX[22][5] ), .Y(n12838) );
  INVX1 U14217 ( .A(\regX[3][5] ), .Y(n12718) );
  OAI22X1 U14218 ( .A(n12867), .B(n14895), .C(n12810), .D(n14896), .Y(n14944)
         );
  INVX1 U14219 ( .A(\regX[24][5] ), .Y(n12810) );
  INVX1 U14220 ( .A(\regX[20][5] ), .Y(n12867) );
  AOI21X1 U14221 ( .A(n14897), .B(\regX[16][5] ), .C(n14946), .Y(n14937) );
  OAI22X1 U14222 ( .A(n13172), .B(n14899), .C(n12877), .D(n14900), .Y(n14946)
         );
  INVX1 U14223 ( .A(\regX[21][5] ), .Y(n12877) );
  OAI21X1 U14224 ( .A(n14947), .B(n13921), .C(n12517), .Y(\U3/U118/Z_4 ) );
  NAND2X1 U14225 ( .A(fGy[4]), .B(n15377), .Y(n12517) );
  NOR2X1 U14226 ( .A(n14948), .B(n14949), .Y(n14947) );
  NAND2X1 U14227 ( .A(n14950), .B(n14951), .Y(n14949) );
  NOR2X1 U14228 ( .A(n14952), .B(n14953), .Y(n14951) );
  OAI21X1 U14229 ( .A(n12674), .B(n14860), .C(n14954), .Y(n14953) );
  AOI22X1 U14230 ( .A(n14862), .B(\regX[11][4] ), .C(n14863), .D(\regX[7][4] ), 
        .Y(n14954) );
  OAI21X1 U14231 ( .A(n12695), .B(n14864), .C(n14955), .Y(n14952) );
  AOI22X1 U14232 ( .A(n14866), .B(N1619), .C(n14867), .D(\regX[23][4] ), .Y(
        n14955) );
  INVX1 U14233 ( .A(\regX[1][4] ), .Y(n12695) );
  NOR2X1 U14234 ( .A(n14956), .B(n14957), .Y(n14950) );
  OAI21X1 U14235 ( .A(n12776), .B(n14870), .C(n14958), .Y(n14957) );
  AOI22X1 U14236 ( .A(n14872), .B(\regX[5][4] ), .C(n14873), .D(\regX[0][4] ), 
        .Y(n14958) );
  INVX1 U14237 ( .A(\regX[9][4] ), .Y(n12776) );
  OAI21X1 U14238 ( .A(n12706), .B(n14874), .C(n14959), .Y(n14956) );
  AOI22X1 U14239 ( .A(n14876), .B(\regX[13][4] ), .C(n14877), .D(N1437), .Y(
        n14959) );
  NAND3X1 U14240 ( .A(n14960), .B(n14961), .C(n14962), .Y(n14948) );
  NOR2X1 U14241 ( .A(n14963), .B(n14964), .Y(n14962) );
  OAI21X1 U14242 ( .A(n12765), .B(n14883), .C(n14965), .Y(n14964) );
  AOI22X1 U14243 ( .A(n14885), .B(N1681), .C(n14886), .D(\regX[17][4] ), .Y(
        n14965) );
  INVX1 U14244 ( .A(\regX[8][4] ), .Y(n12765) );
  OAI21X1 U14245 ( .A(n12585), .B(n14887), .C(n14966), .Y(n14963) );
  AOI22X1 U14246 ( .A(n14889), .B(N1739), .C(n14890), .D(\regX[19][4] ), .Y(
        n14966) );
  INVX1 U14247 ( .A(\regX[15][4] ), .Y(n12585) );
  NOR2X1 U14248 ( .A(n14967), .B(n14968), .Y(n14961) );
  OAI22X1 U14249 ( .A(n12717), .B(n14893), .C(n12837), .D(n14894), .Y(n14968)
         );
  INVX1 U14250 ( .A(\regX[22][4] ), .Y(n12837) );
  INVX1 U14251 ( .A(\regX[3][4] ), .Y(n12717) );
  OAI22X1 U14252 ( .A(n12866), .B(n14895), .C(n12809), .D(n14896), .Y(n14967)
         );
  INVX1 U14253 ( .A(\regX[24][4] ), .Y(n12809) );
  INVX1 U14254 ( .A(\regX[20][4] ), .Y(n12866) );
  AOI21X1 U14255 ( .A(n14897), .B(\regX[16][4] ), .C(n14969), .Y(n14960) );
  OAI22X1 U14256 ( .A(n13171), .B(n14899), .C(n12876), .D(n14900), .Y(n14969)
         );
  INVX1 U14257 ( .A(\regX[21][4] ), .Y(n12876) );
  NOR2X1 U14258 ( .A(n14214), .B(n13030), .Y(\U3/U118/Z_31 ) );
  INVX1 U14259 ( .A(fGy[31]), .Y(n13030) );
  NOR2X1 U14260 ( .A(n14214), .B(n13028), .Y(\U3/U118/Z_30 ) );
  INVX1 U14261 ( .A(fGy[30]), .Y(n13028) );
  OAI21X1 U14262 ( .A(n14214), .B(n14595), .C(n14970), .Y(\U3/U118/Z_3 ) );
  AOI21X1 U14263 ( .A(n15369), .B(n14971), .C(n15328), .Y(n14970) );
  NAND3X1 U14264 ( .A(n14972), .B(n14973), .C(n14974), .Y(n14971) );
  NOR2X1 U14265 ( .A(n14975), .B(n14976), .Y(n14974) );
  OR2X1 U14266 ( .A(n14977), .B(n14978), .Y(n14976) );
  OAI21X1 U14267 ( .A(n12764), .B(n14883), .C(n14979), .Y(n14978) );
  AOI22X1 U14268 ( .A(n14885), .B(N1680), .C(n14886), .D(\regX[17][3] ), .Y(
        n14979) );
  INVX1 U14269 ( .A(\regX[8][3] ), .Y(n12764) );
  OAI21X1 U14270 ( .A(n12583), .B(n14887), .C(n14980), .Y(n14977) );
  AOI22X1 U14271 ( .A(n14889), .B(N1738), .C(n14890), .D(\regX[19][3] ), .Y(
        n14980) );
  INVX1 U14272 ( .A(\regX[15][3] ), .Y(n12583) );
  NAND3X1 U14273 ( .A(n14981), .B(n14982), .C(n14983), .Y(n14975) );
  AOI21X1 U14274 ( .A(n14897), .B(\regX[16][3] ), .C(n14984), .Y(n14983) );
  OAI22X1 U14275 ( .A(n13170), .B(n14899), .C(n12875), .D(n14900), .Y(n14984)
         );
  INVX1 U14276 ( .A(\regX[21][3] ), .Y(n12875) );
  AOI22X1 U14277 ( .A(n14985), .B(\regX[24][3] ), .C(n14986), .D(\regX[20][3] ), .Y(n14982) );
  AOI22X1 U14278 ( .A(n14987), .B(\regX[22][3] ), .C(n14988), .D(\regX[3][3] ), 
        .Y(n14981) );
  NOR2X1 U14279 ( .A(n14989), .B(n14990), .Y(n14973) );
  OAI21X1 U14280 ( .A(n12673), .B(n14860), .C(n14991), .Y(n14990) );
  AOI22X1 U14281 ( .A(n14862), .B(\regX[11][3] ), .C(n14863), .D(\regX[7][3] ), 
        .Y(n14991) );
  OAI21X1 U14282 ( .A(n12694), .B(n14864), .C(n14992), .Y(n14989) );
  AOI22X1 U14283 ( .A(n14866), .B(N1618), .C(n14867), .D(\regX[23][3] ), .Y(
        n14992) );
  INVX1 U14284 ( .A(\regX[1][3] ), .Y(n12694) );
  NOR2X1 U14285 ( .A(n14993), .B(n14994), .Y(n14972) );
  OAI21X1 U14286 ( .A(n12775), .B(n14870), .C(n14995), .Y(n14994) );
  AOI22X1 U14287 ( .A(n14872), .B(\regX[5][3] ), .C(n14873), .D(\regX[0][3] ), 
        .Y(n14995) );
  INVX1 U14288 ( .A(\regX[9][3] ), .Y(n12775) );
  OAI21X1 U14289 ( .A(n12705), .B(n14874), .C(n14996), .Y(n14993) );
  AOI22X1 U14290 ( .A(n14876), .B(\regX[13][3] ), .C(n14877), .D(N1436), .Y(
        n14996) );
  NOR2X1 U14291 ( .A(n14214), .B(n13026), .Y(\U3/U118/Z_29 ) );
  INVX1 U14292 ( .A(fGy[29]), .Y(n13026) );
  NOR2X1 U14293 ( .A(n14214), .B(n13024), .Y(\U3/U118/Z_28 ) );
  INVX1 U14294 ( .A(fGy[28]), .Y(n13024) );
  NOR2X1 U14295 ( .A(n14214), .B(n13022), .Y(\U3/U118/Z_27 ) );
  INVX1 U14296 ( .A(fGy[27]), .Y(n13022) );
  NOR2X1 U14297 ( .A(n14214), .B(n13020), .Y(\U3/U118/Z_26 ) );
  INVX1 U14298 ( .A(fGy[26]), .Y(n13020) );
  NOR2X1 U14299 ( .A(n14214), .B(n13018), .Y(\U3/U118/Z_25 ) );
  INVX1 U14300 ( .A(fGy[25]), .Y(n13018) );
  NOR2X1 U14301 ( .A(n14214), .B(n13016), .Y(\U3/U118/Z_24 ) );
  INVX1 U14302 ( .A(fGy[24]), .Y(n13016) );
  NOR2X1 U14303 ( .A(n14214), .B(n13014), .Y(\U3/U118/Z_23 ) );
  INVX1 U14304 ( .A(fGy[23]), .Y(n13014) );
  NOR2X1 U14305 ( .A(n14214), .B(n13012), .Y(\U3/U118/Z_22 ) );
  INVX1 U14306 ( .A(fGy[22]), .Y(n13012) );
  NOR2X1 U14307 ( .A(n14214), .B(n13010), .Y(\U3/U118/Z_21 ) );
  INVX1 U14308 ( .A(fGy[21]), .Y(n13010) );
  NOR2X1 U14309 ( .A(n14214), .B(n13008), .Y(\U3/U118/Z_20 ) );
  INVX1 U14310 ( .A(fGy[20]), .Y(n13008) );
  NAND3X1 U14311 ( .A(n12552), .B(n14997), .C(n14998), .Y(\U3/U118/Z_2 ) );
  OAI21X1 U14312 ( .A(n14999), .B(n15000), .C(n15369), .Y(n14998) );
  NAND2X1 U14313 ( .A(n15001), .B(n15002), .Y(n15000) );
  NOR2X1 U14314 ( .A(n15003), .B(n15004), .Y(n15002) );
  OAI21X1 U14315 ( .A(n12672), .B(n14860), .C(n15005), .Y(n15004) );
  AOI22X1 U14316 ( .A(n14862), .B(\regX[11][2] ), .C(n14863), .D(\regX[7][2] ), 
        .Y(n15005) );
  OAI21X1 U14317 ( .A(n12693), .B(n14864), .C(n15006), .Y(n15003) );
  AOI22X1 U14318 ( .A(n14866), .B(N1617), .C(n14867), .D(\regX[23][2] ), .Y(
        n15006) );
  INVX1 U14319 ( .A(\regX[1][2] ), .Y(n12693) );
  NOR2X1 U14320 ( .A(n15007), .B(n15008), .Y(n15001) );
  OAI21X1 U14321 ( .A(n12774), .B(n14870), .C(n15009), .Y(n15008) );
  AOI22X1 U14322 ( .A(n14872), .B(\regX[5][2] ), .C(n14873), .D(\regX[0][2] ), 
        .Y(n15009) );
  INVX1 U14323 ( .A(\regX[9][2] ), .Y(n12774) );
  OAI21X1 U14324 ( .A(n12704), .B(n14874), .C(n15010), .Y(n15007) );
  AOI22X1 U14325 ( .A(n14876), .B(\regX[13][2] ), .C(n14877), .D(N1435), .Y(
        n15010) );
  NAND3X1 U14326 ( .A(n15011), .B(n15012), .C(n15013), .Y(n14999) );
  NOR2X1 U14327 ( .A(n15014), .B(n15015), .Y(n15013) );
  OAI21X1 U14328 ( .A(n12763), .B(n14883), .C(n15016), .Y(n15015) );
  AOI22X1 U14329 ( .A(n14885), .B(N1679), .C(n14886), .D(\regX[17][2] ), .Y(
        n15016) );
  INVX1 U14330 ( .A(\regX[8][2] ), .Y(n12763) );
  OAI21X1 U14331 ( .A(n12581), .B(n14887), .C(n15017), .Y(n15014) );
  AOI22X1 U14332 ( .A(n14889), .B(N1737), .C(n14890), .D(\regX[19][2] ), .Y(
        n15017) );
  INVX1 U14333 ( .A(\regX[15][2] ), .Y(n12581) );
  NOR2X1 U14334 ( .A(n15018), .B(n15019), .Y(n15012) );
  OAI22X1 U14335 ( .A(n12715), .B(n14893), .C(n12835), .D(n14894), .Y(n15019)
         );
  INVX1 U14336 ( .A(\regX[22][2] ), .Y(n12835) );
  INVX1 U14337 ( .A(\regX[3][2] ), .Y(n12715) );
  OAI22X1 U14338 ( .A(n12864), .B(n14895), .C(n12807), .D(n14896), .Y(n15018)
         );
  INVX1 U14339 ( .A(\regX[24][2] ), .Y(n12807) );
  INVX1 U14340 ( .A(\regX[20][2] ), .Y(n12864) );
  AOI21X1 U14341 ( .A(n14897), .B(\regX[16][2] ), .C(n15020), .Y(n15011) );
  OAI22X1 U14342 ( .A(n13169), .B(n14899), .C(n12874), .D(n14900), .Y(n15020)
         );
  INVX1 U14343 ( .A(\regX[21][2] ), .Y(n12874) );
  INVX1 U14344 ( .A(n15375), .Y(n14997) );
  NOR2X1 U14345 ( .A(n14596), .B(n14214), .Y(n15375) );
  INVX1 U14346 ( .A(fGy[2]), .Y(n14596) );
  NOR2X1 U14347 ( .A(n14214), .B(n13006), .Y(\U3/U118/Z_19 ) );
  INVX1 U14348 ( .A(fGy[19]), .Y(n13006) );
  NOR2X1 U14349 ( .A(n14214), .B(n13004), .Y(\U3/U118/Z_18 ) );
  INVX1 U14350 ( .A(fGy[18]), .Y(n13004) );
  NOR2X1 U14351 ( .A(n14214), .B(n13002), .Y(\U3/U118/Z_17 ) );
  INVX1 U14352 ( .A(fGy[17]), .Y(n13002) );
  NOR2X1 U14353 ( .A(n14214), .B(n13000), .Y(\U3/U118/Z_16 ) );
  INVX1 U14354 ( .A(fGy[16]), .Y(n13000) );
  NOR2X1 U14355 ( .A(n14214), .B(n12998), .Y(\U3/U118/Z_15 ) );
  INVX1 U14356 ( .A(fGy[15]), .Y(n12998) );
  NOR2X1 U14357 ( .A(n14214), .B(n12996), .Y(\U3/U118/Z_14 ) );
  INVX1 U14358 ( .A(fGy[14]), .Y(n12996) );
  NOR2X1 U14359 ( .A(n14214), .B(n12994), .Y(\U3/U118/Z_13 ) );
  INVX1 U14360 ( .A(fGy[13]), .Y(n12994) );
  NOR2X1 U14361 ( .A(n14214), .B(n12992), .Y(\U3/U118/Z_12 ) );
  INVX1 U14362 ( .A(fGy[12]), .Y(n12992) );
  NOR2X1 U14363 ( .A(n14214), .B(n12990), .Y(\U3/U118/Z_11 ) );
  INVX1 U14364 ( .A(fGy[11]), .Y(n12990) );
  NOR2X1 U14365 ( .A(n14214), .B(n12988), .Y(\U3/U118/Z_10 ) );
  INVX1 U14366 ( .A(fGy[10]), .Y(n12988) );
  OAI21X1 U14367 ( .A(n14214), .B(n14597), .C(n15021), .Y(\U3/U118/Z_1 ) );
  AOI21X1 U14368 ( .A(n15369), .B(n15022), .C(n15328), .Y(n15021) );
  NAND3X1 U14369 ( .A(n15023), .B(n15024), .C(n15025), .Y(n15022) );
  NOR2X1 U14370 ( .A(n15026), .B(n15027), .Y(n15025) );
  OR2X1 U14371 ( .A(n15028), .B(n15029), .Y(n15027) );
  OAI21X1 U14372 ( .A(n12762), .B(n14883), .C(n15030), .Y(n15029) );
  AOI22X1 U14373 ( .A(n14885), .B(N1678), .C(n14886), .D(\regX[17][1] ), .Y(
        n15030) );
  INVX1 U14374 ( .A(\regX[8][1] ), .Y(n12762) );
  OAI21X1 U14375 ( .A(n12579), .B(n14887), .C(n15031), .Y(n15028) );
  AOI22X1 U14376 ( .A(n14889), .B(N1736), .C(n14890), .D(\regX[19][1] ), .Y(
        n15031) );
  INVX1 U14377 ( .A(\regX[15][1] ), .Y(n12579) );
  NAND3X1 U14378 ( .A(n15032), .B(n15033), .C(n15034), .Y(n15026) );
  AOI21X1 U14379 ( .A(n14897), .B(\regX[16][1] ), .C(n15035), .Y(n15034) );
  OAI22X1 U14380 ( .A(n13168), .B(n14899), .C(n12873), .D(n14900), .Y(n15035)
         );
  INVX1 U14381 ( .A(\regX[21][1] ), .Y(n12873) );
  AOI22X1 U14382 ( .A(n14985), .B(\regX[24][1] ), .C(n14986), .D(\regX[20][1] ), .Y(n15033) );
  INVX1 U14383 ( .A(n14895), .Y(n14986) );
  AOI22X1 U14384 ( .A(n14987), .B(\regX[22][1] ), .C(n14988), .D(\regX[3][1] ), 
        .Y(n15032) );
  INVX1 U14385 ( .A(n14893), .Y(n14988) );
  INVX1 U14386 ( .A(n14894), .Y(n14987) );
  NOR2X1 U14387 ( .A(n15036), .B(n15037), .Y(n15024) );
  OAI21X1 U14388 ( .A(n12671), .B(n14860), .C(n15038), .Y(n15037) );
  AOI22X1 U14389 ( .A(n14862), .B(\regX[11][1] ), .C(n14863), .D(\regX[7][1] ), 
        .Y(n15038) );
  OAI21X1 U14390 ( .A(n12692), .B(n14864), .C(n15039), .Y(n15036) );
  AOI22X1 U14391 ( .A(n14866), .B(N1616), .C(n14867), .D(\regX[23][1] ), .Y(
        n15039) );
  INVX1 U14392 ( .A(\regX[1][1] ), .Y(n12692) );
  NOR2X1 U14393 ( .A(n15040), .B(n15041), .Y(n15023) );
  OAI21X1 U14394 ( .A(n12773), .B(n14870), .C(n15042), .Y(n15041) );
  AOI22X1 U14395 ( .A(n14872), .B(\regX[5][1] ), .C(n14873), .D(\regX[0][1] ), 
        .Y(n15042) );
  INVX1 U14396 ( .A(\regX[9][1] ), .Y(n12773) );
  OAI21X1 U14397 ( .A(n12703), .B(n14874), .C(n15043), .Y(n15040) );
  AOI22X1 U14398 ( .A(n14876), .B(\regX[13][1] ), .C(n14877), .D(N1434), .Y(
        n15043) );
  NAND3X1 U14399 ( .A(n12552), .B(n15044), .C(n15045), .Y(\U3/U118/Z_0 ) );
  OAI21X1 U14400 ( .A(n15046), .B(n15047), .C(n15369), .Y(n15045) );
  NAND2X1 U14401 ( .A(n15048), .B(n15049), .Y(n15047) );
  NOR2X1 U14402 ( .A(n15050), .B(n15051), .Y(n15049) );
  OAI21X1 U14403 ( .A(n12669), .B(n14860), .C(n15052), .Y(n15051) );
  AOI22X1 U14404 ( .A(n14862), .B(\regX[11][0] ), .C(n14863), .D(\regX[7][0] ), 
        .Y(n15052) );
  AND2X1 U14405 ( .A(n15053), .B(n15054), .Y(n14863) );
  AND2X1 U14406 ( .A(n15055), .B(n15056), .Y(n14862) );
  NAND2X1 U14407 ( .A(n15057), .B(n15054), .Y(n14860) );
  OAI21X1 U14408 ( .A(n12690), .B(n14864), .C(n15058), .Y(n15050) );
  AOI22X1 U14409 ( .A(n14866), .B(N1615), .C(n14867), .D(\regX[23][0] ), .Y(
        n15058) );
  AND2X1 U14410 ( .A(n15059), .B(n15054), .Y(n14867) );
  AND2X1 U14411 ( .A(n15060), .B(n15056), .Y(n14866) );
  NAND2X1 U14412 ( .A(n15061), .B(n15053), .Y(n14864) );
  INVX1 U14413 ( .A(\regX[1][0] ), .Y(n12690) );
  NOR2X1 U14414 ( .A(n15062), .B(n15063), .Y(n15048) );
  OAI21X1 U14415 ( .A(n12771), .B(n14870), .C(n15064), .Y(n15063) );
  AOI22X1 U14416 ( .A(n14872), .B(\regX[5][0] ), .C(n14873), .D(\regX[0][0] ), 
        .Y(n15064) );
  AND2X1 U14417 ( .A(n15057), .B(n15061), .Y(n14873) );
  AND2X1 U14418 ( .A(n15053), .B(n15065), .Y(n14872) );
  NAND2X1 U14419 ( .A(n15055), .B(n15061), .Y(n14870) );
  INVX1 U14420 ( .A(\regX[9][0] ), .Y(n12771) );
  OAI21X1 U14421 ( .A(n12701), .B(n14874), .C(n15066), .Y(n15062) );
  AOI22X1 U14422 ( .A(n14876), .B(\regX[13][0] ), .C(n14877), .D(N1433), .Y(
        n15066) );
  AND2X1 U14423 ( .A(n15057), .B(n15065), .Y(n14877) );
  AND2X1 U14424 ( .A(n15055), .B(n15065), .Y(n14876) );
  NAND2X1 U14425 ( .A(n15057), .B(n15056), .Y(n14874) );
  INVX1 U14426 ( .A(n15067), .Y(n15057) );
  NAND3X1 U14427 ( .A(n15068), .B(n15069), .C(n15070), .Y(n15067) );
  NAND3X1 U14428 ( .A(n15071), .B(n15072), .C(n15073), .Y(n15046) );
  NOR2X1 U14429 ( .A(n15074), .B(n15075), .Y(n15073) );
  OAI21X1 U14430 ( .A(n12760), .B(n14883), .C(n15076), .Y(n15075) );
  AOI22X1 U14431 ( .A(n14885), .B(N1677), .C(n14886), .D(\regX[17][0] ), .Y(
        n15076) );
  AND2X1 U14432 ( .A(n15061), .B(n15059), .Y(n14886) );
  AND2X1 U14433 ( .A(n15060), .B(n15065), .Y(n14885) );
  NAND3X1 U14434 ( .A(n15061), .B(n15068), .C(n15060), .Y(n14883) );
  INVX1 U14435 ( .A(\regX[8][0] ), .Y(n12760) );
  OAI21X1 U14436 ( .A(n12576), .B(n14887), .C(n15077), .Y(n15074) );
  AOI22X1 U14437 ( .A(n14889), .B(N1735), .C(n14890), .D(\regX[19][0] ), .Y(
        n15077) );
  AND2X1 U14438 ( .A(n15059), .B(n15056), .Y(n14890) );
  AND2X1 U14439 ( .A(n15060), .B(n15054), .Y(n14889) );
  NOR2X1 U14440 ( .A(n15078), .B(n15069), .Y(n15060) );
  NAND2X1 U14441 ( .A(n15055), .B(n15054), .Y(n14887) );
  NOR2X1 U14442 ( .A(n15069), .B(n15070), .Y(n15055) );
  INVX1 U14443 ( .A(\regX[15][0] ), .Y(n12576) );
  NOR2X1 U14444 ( .A(n15079), .B(n15080), .Y(n15072) );
  OAI22X1 U14445 ( .A(n12712), .B(n14893), .C(n12832), .D(n14894), .Y(n15080)
         );
  NAND2X1 U14446 ( .A(n15054), .B(n15081), .Y(n14894) );
  NOR2X1 U14447 ( .A(n15082), .B(n15083), .Y(n15054) );
  INVX1 U14448 ( .A(\regX[22][0] ), .Y(n12832) );
  NAND2X1 U14449 ( .A(n15056), .B(n15053), .Y(n14893) );
  INVX1 U14450 ( .A(n15084), .Y(n15053) );
  NAND3X1 U14451 ( .A(n15068), .B(n15069), .C(n15078), .Y(n15084) );
  INVX1 U14452 ( .A(\regX[3][0] ), .Y(n12712) );
  OAI22X1 U14453 ( .A(n12861), .B(n14895), .C(n12804), .D(n14896), .Y(n15079)
         );
  INVX1 U14454 ( .A(n14985), .Y(n14896) );
  NOR2X1 U14455 ( .A(n15069), .B(n15068), .Y(n14985) );
  INVX1 U14456 ( .A(\regX[24][0] ), .Y(n12804) );
  NAND2X1 U14457 ( .A(n15065), .B(n15081), .Y(n14895) );
  INVX1 U14458 ( .A(\regX[20][0] ), .Y(n12861) );
  AOI21X1 U14459 ( .A(n14897), .B(\regX[16][0] ), .C(n15085), .Y(n15071) );
  OAI22X1 U14460 ( .A(n12555), .B(n14899), .C(n12871), .D(n14900), .Y(n15085)
         );
  NAND2X1 U14461 ( .A(n15059), .B(n15065), .Y(n14900) );
  NOR2X1 U14462 ( .A(n15086), .B(n15083), .Y(n15065) );
  NOR2X1 U14463 ( .A(n15068), .B(n15070), .Y(n15059) );
  INVX1 U14464 ( .A(n15078), .Y(n15070) );
  INVX1 U14465 ( .A(\regX[21][0] ), .Y(n12871) );
  NAND2X1 U14466 ( .A(n15056), .B(n15081), .Y(n14899) );
  NOR2X1 U14467 ( .A(n15087), .B(n15082), .Y(n15056) );
  INVX1 U14468 ( .A(\regX[18][0] ), .Y(n12555) );
  INVX1 U14469 ( .A(n15088), .Y(n14897) );
  NAND3X1 U14470 ( .A(n15081), .B(n15069), .C(n15061), .Y(n15088) );
  NOR2X1 U14471 ( .A(n15087), .B(n15086), .Y(n15061) );
  INVX1 U14472 ( .A(n15082), .Y(n15086) );
  XOR2X1 U14473 ( .A(n15089), .B(n14569), .Y(n15082) );
  INVX1 U14474 ( .A(n14572), .Y(n14569) );
  NAND2X1 U14475 ( .A(n15090), .B(n15091), .Y(n15089) );
  OAI21X1 U14476 ( .A(n14563), .B(n15092), .C(n15093), .Y(n15091) );
  INVX1 U14477 ( .A(N3090), .Y(n15093) );
  INVX1 U14478 ( .A(n15083), .Y(n15087) );
  AOI21X1 U14479 ( .A(n15094), .B(N3091), .C(n15095), .Y(n15083) );
  XNOR2X1 U14480 ( .A(N3092), .B(n15096), .Y(n15069) );
  NOR2X1 U14481 ( .A(n15078), .B(n15068), .Y(n15081) );
  XNOR2X1 U14482 ( .A(n15097), .B(N3093), .Y(n15068) );
  OAI21X1 U14483 ( .A(n15095), .B(n14562), .C(n15098), .Y(n15097) );
  OAI21X1 U14484 ( .A(n15099), .B(n15096), .C(N3092), .Y(n15098) );
  INVX1 U14485 ( .A(n15095), .Y(n15096) );
  INVX1 U14486 ( .A(n14562), .Y(n15099) );
  XNOR2X1 U14487 ( .A(n15100), .B(n14578), .Y(n14562) );
  XNOR2X1 U14488 ( .A(n14591), .B(n14588), .Y(n15100) );
  INVX1 U14489 ( .A(n14592), .Y(n14588) );
  OAI21X1 U14490 ( .A(n14594), .B(n14193), .C(n15101), .Y(n14592) );
  OAI21X1 U14491 ( .A(n14200), .B(n15102), .C(n14578), .Y(n15101) );
  INVX1 U14492 ( .A(n14200), .Y(n14193) );
  XOR2X1 U14493 ( .A(n15103), .B(n15104), .Y(n14200) );
  XNOR2X1 U14494 ( .A(n15105), .B(n15106), .Y(n15104) );
  INVX1 U14495 ( .A(n15102), .Y(n14594) );
  OAI21X1 U14496 ( .A(n15107), .B(n15108), .C(n15109), .Y(n15102) );
  OAI21X1 U14497 ( .A(n15110), .B(n15111), .C(n14578), .Y(n15109) );
  INVX1 U14498 ( .A(n15107), .Y(n15111) );
  NOR2X1 U14499 ( .A(n14170), .B(n12552), .Y(n14591) );
  XOR2X1 U14500 ( .A(n15112), .B(n14587), .Y(n14170) );
  OAI21X1 U14501 ( .A(n15103), .B(n15113), .C(n15114), .Y(n14587) );
  OAI21X1 U14502 ( .A(n15105), .B(n15115), .C(n15106), .Y(n15114) );
  OAI21X1 U14503 ( .A(n15116), .B(n15117), .C(n15118), .Y(n15106) );
  OAI21X1 U14504 ( .A(n15119), .B(n15120), .C(n15121), .Y(n15118) );
  INVX1 U14505 ( .A(n15116), .Y(n15120) );
  INVX1 U14506 ( .A(n15119), .Y(n15117) );
  INVX1 U14507 ( .A(n15103), .Y(n15115) );
  INVX1 U14508 ( .A(n15113), .Y(n15105) );
  OAI21X1 U14509 ( .A(n13921), .B(n15122), .C(n15123), .Y(n15113) );
  INVX1 U14510 ( .A(N3091), .Y(n15122) );
  NOR2X1 U14511 ( .A(n14828), .B(n15328), .Y(n15103) );
  XOR2X1 U14512 ( .A(n15124), .B(n15125), .Y(n14828) );
  XNOR2X1 U14513 ( .A(n15126), .B(n15127), .Y(n15124) );
  OAI21X1 U14514 ( .A(n14585), .B(n14586), .C(n14584), .Y(n15112) );
  NAND2X1 U14515 ( .A(n14585), .B(n14586), .Y(n14584) );
  NOR2X1 U14516 ( .A(n14809), .B(n13921), .Y(n14586) );
  XOR2X1 U14517 ( .A(n15128), .B(n14849), .Y(n14809) );
  MUX2X1 U14518 ( .B(n15129), .A(n14847), .S(n14845), .Y(n14849) );
  NOR2X1 U14519 ( .A(N3342), .B(n12552), .Y(n15129) );
  XNOR2X1 U14520 ( .A(n14838), .B(n14848), .Y(n15128) );
  INVX1 U14521 ( .A(n14851), .Y(n14848) );
  OAI21X1 U14522 ( .A(n15126), .B(n15127), .C(n15130), .Y(n14851) );
  OAI21X1 U14523 ( .A(n15131), .B(n15132), .C(n14838), .Y(n15130) );
  INVX1 U14524 ( .A(n15132), .Y(n15127) );
  OAI21X1 U14525 ( .A(n15133), .B(n15123), .C(n15134), .Y(n15132) );
  NOR2X1 U14526 ( .A(n14845), .B(n15369), .Y(n15134) );
  NOR2X1 U14527 ( .A(N3340), .B(N3341), .Y(n14845) );
  NAND2X1 U14528 ( .A(N3341), .B(n15328), .Y(n15123) );
  INVX1 U14529 ( .A(n15131), .Y(n15126) );
  OAI21X1 U14530 ( .A(n15135), .B(n15125), .C(n15136), .Y(n15131) );
  OAI21X1 U14531 ( .A(n14838), .B(n15137), .C(n15138), .Y(n15136) );
  INVX1 U14532 ( .A(n15135), .Y(n15137) );
  INVX1 U14533 ( .A(n14838), .Y(n15125) );
  AOI21X1 U14534 ( .A(n15369), .B(N3092), .C(n14847), .Y(n14585) );
  NOR2X1 U14535 ( .A(n14846), .B(n12552), .Y(n14847) );
  INVX1 U14536 ( .A(N3342), .Y(n14846) );
  NOR2X1 U14537 ( .A(n15094), .B(N3091), .Y(n15095) );
  OAI21X1 U14538 ( .A(n15139), .B(n14572), .C(n15090), .Y(n15094) );
  NAND3X1 U14539 ( .A(N3090), .B(n14565), .C(N3089), .Y(n15090) );
  XNOR2X1 U14540 ( .A(n15140), .B(n14578), .Y(n14572) );
  XNOR2X1 U14541 ( .A(n12552), .B(dx[1]), .Y(n14578) );
  XNOR2X1 U14542 ( .A(n15110), .B(n15107), .Y(n15140) );
  NOR2X1 U14543 ( .A(n14199), .B(n15369), .Y(n15107) );
  XOR2X1 U14544 ( .A(n15119), .B(n15141), .Y(n14199) );
  XNOR2X1 U14545 ( .A(n15116), .B(n15121), .Y(n15141) );
  NOR2X1 U14546 ( .A(n14829), .B(n15328), .Y(n15116) );
  XOR2X1 U14547 ( .A(n15142), .B(n15138), .Y(n14829) );
  XNOR2X1 U14548 ( .A(n14838), .B(n15135), .Y(n15142) );
  NOR2X1 U14549 ( .A(n15133), .B(n15369), .Y(n15135) );
  INVX1 U14550 ( .A(N3340), .Y(n15133) );
  XNOR2X1 U14551 ( .A(dx[1]), .B(n13921), .Y(n14838) );
  AOI22X1 U14552 ( .A(n15328), .B(N3340), .C(n15369), .D(N3090), .Y(n15119) );
  INVX1 U14553 ( .A(n15108), .Y(n15110) );
  OAI21X1 U14554 ( .A(n14186), .B(n15143), .C(n15328), .Y(n15108) );
  AOI21X1 U14555 ( .A(N3089), .B(n14565), .C(N3090), .Y(n15139) );
  XNOR2X1 U14556 ( .A(N3089), .B(n14563), .Y(n15078) );
  INVX1 U14557 ( .A(n14565), .Y(n14563) );
  XOR2X1 U14558 ( .A(n15143), .B(n15144), .Y(n14565) );
  NOR2X1 U14559 ( .A(n12552), .B(n14186), .Y(n15144) );
  OAI21X1 U14560 ( .A(n15145), .B(n15146), .C(n15121), .Y(n14186) );
  OAI21X1 U14561 ( .A(n13921), .B(n14826), .C(n15145), .Y(n15121) );
  INVX1 U14562 ( .A(n14818), .Y(n14826) );
  NAND2X1 U14563 ( .A(n14818), .B(n15369), .Y(n15146) );
  AOI21X1 U14564 ( .A(n13634), .B(n15147), .C(n15138), .Y(n14818) );
  MUX2X1 U14565 ( .B(dx[0]), .A(n15148), .S(n13921), .Y(n15138) );
  NAND2X1 U14566 ( .A(N3359), .B(dx[0]), .Y(n15148) );
  OAI22X1 U14567 ( .A(n12552), .B(n15147), .C(n13921), .D(n15092), .Y(n15145)
         );
  INVX1 U14568 ( .A(N3089), .Y(n15092) );
  INVX1 U14569 ( .A(N3359), .Y(n15147) );
  XNOR2X1 U14570 ( .A(n15328), .B(n13634), .Y(n15143) );
  INVX1 U14571 ( .A(n15376), .Y(n15044) );
  NOR2X1 U14572 ( .A(n14598), .B(n14214), .Y(n15376) );
  INVX1 U14573 ( .A(fGy[0]), .Y(n14598) );
  OAI21X1 U14574 ( .A(n12470), .B(n13174), .C(n15149), .Y(\U3/U110/Z_7 ) );
  INVX1 U14575 ( .A(\regX[18][7] ), .Y(n13174) );
  OAI21X1 U14576 ( .A(n12470), .B(n13173), .C(n15149), .Y(\U3/U110/Z_6 ) );
  INVX1 U14577 ( .A(\regX[18][6] ), .Y(n13173) );
  OAI21X1 U14578 ( .A(n12470), .B(n13172), .C(n15149), .Y(\U3/U110/Z_5 ) );
  INVX1 U14579 ( .A(\regX[18][5] ), .Y(n13172) );
  OAI21X1 U14580 ( .A(n12470), .B(n13171), .C(n15149), .Y(\U3/U110/Z_4 ) );
  INVX1 U14581 ( .A(\regX[18][4] ), .Y(n13171) );
  OAI21X1 U14582 ( .A(n12470), .B(n13170), .C(n15149), .Y(\U3/U110/Z_3 ) );
  INVX1 U14583 ( .A(\regX[18][3] ), .Y(n13170) );
  OAI21X1 U14584 ( .A(n12470), .B(n13169), .C(n15149), .Y(\U3/U110/Z_2 ) );
  INVX1 U14585 ( .A(\regX[18][2] ), .Y(n13169) );
  OAI21X1 U14586 ( .A(n12470), .B(n13168), .C(n15149), .Y(\U3/U110/Z_1 ) );
  NAND2X1 U14587 ( .A(dy[1]), .B(n15328), .Y(n15149) );
  INVX1 U14588 ( .A(\regX[18][1] ), .Y(n13168) );
  NAND2X1 U14589 ( .A(n12552), .B(n12470), .Y(\U3/U109/Z_2 ) );
  NAND3X1 U14590 ( .A(n13653), .B(n12646), .C(n12471), .Y(n12554) );
  INVX1 U14591 ( .A(n15328), .Y(n12552) );
  OAI21X1 U14592 ( .A(n14214), .B(n14595), .C(n15150), .Y(\U3/U106/Z_3 ) );
  INVX1 U14593 ( .A(fGy[3]), .Y(n14595) );
  OAI21X1 U14594 ( .A(n14214), .B(n14597), .C(n15150), .Y(\U3/U106/Z_1 ) );
  INVX1 U14595 ( .A(fGy[1]), .Y(n14597) );
  OAI22X1 U14596 ( .A(n12673), .B(n15150), .C(n14214), .D(n14295), .Y(
        \U3/U105/Z_3 ) );
  INVX1 U14597 ( .A(N2749), .Y(n14295) );
  INVX1 U14598 ( .A(\regX[6][3] ), .Y(n12673) );
  OAI22X1 U14599 ( .A(n12672), .B(n15150), .C(n14214), .D(n14297), .Y(
        \U3/U105/Z_2 ) );
  INVX1 U14600 ( .A(N2748), .Y(n14297) );
  INVX1 U14601 ( .A(\regX[6][2] ), .Y(n12672) );
  OAI22X1 U14602 ( .A(n12671), .B(n15150), .C(n14214), .D(n14308), .Y(
        \U3/U105/Z_1 ) );
  INVX1 U14603 ( .A(N2747), .Y(n14308) );
  INVX1 U14604 ( .A(\regX[6][1] ), .Y(n12671) );
  OAI22X1 U14605 ( .A(n12669), .B(n15150), .C(n14214), .D(n14319), .Y(
        \U3/U105/Z_0 ) );
  INVX1 U14606 ( .A(N2746), .Y(n14319) );
  INVX1 U14607 ( .A(\regX[6][0] ), .Y(n12669) );
  NOR2X1 U14608 ( .A(n12556), .B(n13399), .Y(\U3/U101/Z_6 ) );
  XOR2X1 U14609 ( .A(n15151), .B(n13590), .Y(n13399) );
  OAI21X1 U14610 ( .A(n13419), .B(n15152), .C(n15153), .Y(n13590) );
  INVX1 U14611 ( .A(N3443), .Y(n15152) );
  XNOR2X1 U14612 ( .A(n15325), .B(n15154), .Y(n15151) );
  NOR2X1 U14613 ( .A(n15155), .B(n15156), .Y(n15154) );
  NOR2X1 U14614 ( .A(n13422), .B(n12556), .Y(\U3/U101/Z_3 ) );
  XNOR2X1 U14615 ( .A(n15156), .B(n15155), .Y(n13422) );
  INVX1 U14616 ( .A(n15157), .Y(n15155) );
  XOR2X1 U14617 ( .A(n13602), .B(n13419), .Y(n15156) );
  OAI21X1 U14618 ( .A(n13419), .B(n15158), .C(n15153), .Y(n13602) );
  INVX1 U14619 ( .A(N3442), .Y(n15158) );
  INVX1 U14620 ( .A(n15159), .Y(\U3/U101/Z_2 ) );
  MUX2X1 U14621 ( .B(n13411), .A(dAddrRegCol[2]), .S(n12556), .Y(n15159) );
  OAI21X1 U14622 ( .A(n15160), .B(n15161), .C(n15157), .Y(n13411) );
  NAND2X1 U14623 ( .A(n15160), .B(n15161), .Y(n15157) );
  XNOR2X1 U14624 ( .A(n13636), .B(n15325), .Y(n15161) );
  OAI21X1 U14625 ( .A(n13419), .B(n15162), .C(n15153), .Y(n13636) );
  MUX2X1 U14626 ( .B(n13418), .A(n15163), .S(n12556), .Y(\U3/U101/Z_1 ) );
  INVX1 U14627 ( .A(dAddrRegCol[1]), .Y(n15163) );
  AOI21X1 U14628 ( .A(n13631), .B(n13632), .C(n15160), .Y(n13418) );
  MUX2X1 U14629 ( .B(n13637), .A(n13638), .S(n13419), .Y(n15160) );
  NAND2X1 U14630 ( .A(n13388), .B(n13638), .Y(n13637) );
  INVX1 U14631 ( .A(n13638), .Y(n13632) );
  OAI21X1 U14632 ( .A(n13419), .B(n15164), .C(n15153), .Y(n13638) );
  NAND2X1 U14633 ( .A(n15327), .B(dx[1]), .Y(n15153) );
  INVX1 U14634 ( .A(n13405), .Y(n15327) );
  INVX1 U14635 ( .A(N1389), .Y(n15164) );
  INVX1 U14636 ( .A(n13388), .Y(n13631) );
  INVX1 U14637 ( .A(n15165), .Y(\U3/U101/Z_0 ) );
  MUX2X1 U14638 ( .B(n13388), .A(dAddrRegCol[0]), .S(n12556), .Y(n15165) );
  OAI21X1 U14639 ( .A(n13405), .B(n13634), .C(n15166), .Y(n13388) );
  NAND2X1 U14640 ( .A(N1388), .B(n15325), .Y(n15166) );
  INVX1 U14641 ( .A(n13419), .Y(n15325) );
  NAND3X1 U14642 ( .A(n15328), .B(n15167), .C(N2880), .Y(n13419) );
  INVX1 U14643 ( .A(N2777), .Y(n15167) );
  NOR2X1 U14644 ( .A(n15150), .B(N3336), .Y(n15328) );
  INVX1 U14645 ( .A(\U3/U107/Z_0 ), .Y(n15150) );
  NOR2X1 U14646 ( .A(n13289), .B(n13165), .Y(\U3/U107/Z_0 ) );
  INVX1 U14647 ( .A(n13058), .Y(n13165) );
  OAI21X1 U14648 ( .A(n14214), .B(n13163), .C(n15168), .Y(n13058) );
  AOI22X1 U14649 ( .A(n15169), .B(n15170), .C(Gy[31]), .D(n12512), .Y(n15168)
         );
  NAND2X1 U14650 ( .A(n12474), .B(n12568), .Y(n12512) );
  NAND3X1 U14651 ( .A(n13166), .B(n12565), .C(IntSignal[1]), .Y(n12568) );
  NAND2X1 U14652 ( .A(n13166), .B(n12537), .Y(n13919) );
  INVX1 U14653 ( .A(n12570), .Y(n13166) );
  NOR2X1 U14654 ( .A(\regX[6][5] ), .B(n15171), .Y(n15170) );
  NAND2X1 U14655 ( .A(n12676), .B(n12677), .Y(n15171) );
  INVX1 U14656 ( .A(\regX[6][7] ), .Y(n12677) );
  INVX1 U14657 ( .A(\regX[6][6] ), .Y(n12676) );
  NOR2X1 U14658 ( .A(n13289), .B(n15172), .Y(n15169) );
  OAI21X1 U14659 ( .A(n15173), .B(n15174), .C(n12674), .Y(n15172) );
  INVX1 U14660 ( .A(\regX[6][4] ), .Y(n12674) );
  NAND2X1 U14661 ( .A(\regX[6][3] ), .B(\regX[6][2] ), .Y(n15174) );
  NAND2X1 U14662 ( .A(\regX[6][1] ), .B(\regX[6][0] ), .Y(n15173) );
  INVX1 U14663 ( .A(fGx[31]), .Y(n13163) );
  NOR2X1 U14664 ( .A(n13892), .B(n12570), .Y(n15377) );
  NAND2X1 U14665 ( .A(n13653), .B(OPMode[0]), .Y(n12570) );
  NOR2X1 U14666 ( .A(OPMode[2]), .B(OPMode[1]), .Y(n13653) );
  NOR2X1 U14667 ( .A(n12510), .B(n12565), .Y(n13911) );
  INVX1 U14668 ( .A(IntSignal[1]), .Y(n12510) );
  NAND3X1 U14669 ( .A(n12537), .B(n12667), .C(OPMode[0]), .Y(n13289) );
  INVX1 U14670 ( .A(dx[0]), .Y(n13634) );
  NAND3X1 U14671 ( .A(n15369), .B(n12687), .C(N2777), .Y(n13405) );
  INVX1 U14672 ( .A(N2549), .Y(n12687) );
  INVX1 U14673 ( .A(n13921), .Y(n15369) );
  NAND3X1 U14674 ( .A(n12667), .B(n12646), .C(n12537), .Y(n13921) );
  NOR2X1 U14675 ( .A(n12565), .B(IntSignal[1]), .Y(n12537) );
  INVX1 U14676 ( .A(IntSignal[0]), .Y(n12565) );
  INVX1 U14677 ( .A(OPMode[0]), .Y(n12646) );
  NOR2X1 U14678 ( .A(n15175), .B(OPMode[2]), .Y(n12667) );
  INVX1 U14679 ( .A(OPMode[1]), .Y(n15175) );
  AND2X1 U14680 ( .A(bCE), .B(N3194), .Y(\U3/U100/Z_6 ) );
  INVX1 U14681 ( .A(n15176), .Y(\U3/U100/Z_4 ) );
  MUX2X1 U14682 ( .B(N3193), .A(N975), .S(n12556), .Y(n15176) );
  INVX1 U14683 ( .A(n15177), .Y(\U3/U100/Z_3 ) );
  MUX2X1 U14684 ( .B(N3192), .A(N974), .S(n12556), .Y(n15177) );
  INVX1 U14685 ( .A(n15178), .Y(\U3/U100/Z_2 ) );
  MUX2X1 U14686 ( .B(N3191), .A(N973), .S(n12556), .Y(n15178) );
  INVX1 U14687 ( .A(n15179), .Y(\U3/U100/Z_1 ) );
  MUX2X1 U14688 ( .B(N3190), .A(N972), .S(n12556), .Y(n15179) );
  INVX1 U14689 ( .A(n15180), .Y(\U3/U100/Z_0 ) );
  MUX2X1 U14690 ( .B(N3189), .A(N971), .S(n12556), .Y(n15180) );
  INVX1 U14691 ( .A(bCE), .Y(n12556) );
  NOR2X1 U14692 ( .A(n15181), .B(n15182), .Y(N1582) );
  OR2X1 U14693 ( .A(n15183), .B(n15184), .Y(n15182) );
  XNOR2X1 U14694 ( .A(n15181), .B(n15185), .Y(N1581) );
  NOR2X1 U14695 ( .A(n15184), .B(n15183), .Y(n15185) );
  INVX1 U14696 ( .A(N1775), .Y(n15183) );
  INVX1 U14697 ( .A(N1776), .Y(n15181) );
  XNOR2X1 U14698 ( .A(N1775), .B(n15184), .Y(N1580) );
  NAND3X1 U14699 ( .A(N1773), .B(n15186), .C(N1774), .Y(n15184) );
  XNOR2X1 U14700 ( .A(N1774), .B(n15187), .Y(N1579) );
  NAND2X1 U14701 ( .A(N1773), .B(n15186), .Y(n15187) );
  XOR2X1 U14702 ( .A(n15186), .B(N1773), .Y(N1578) );
  OAI21X1 U14703 ( .A(n15188), .B(n12829), .C(n15189), .Y(n15186) );
  OAI21X1 U14704 ( .A(N1742), .B(n15190), .C(N1772), .Y(n15189) );
  XNOR2X1 U14705 ( .A(n15188), .B(n15191), .Y(N1577) );
  XNOR2X1 U14706 ( .A(N1772), .B(n12829), .Y(n15191) );
  INVX1 U14707 ( .A(N1742), .Y(n12829) );
  INVX1 U14708 ( .A(n15190), .Y(n15188) );
  OAI21X1 U14709 ( .A(n15192), .B(n12828), .C(n15193), .Y(n15190) );
  OAI21X1 U14710 ( .A(N1741), .B(n15194), .C(N1771), .Y(n15193) );
  INVX1 U14711 ( .A(N1741), .Y(n12828) );
  INVX1 U14712 ( .A(n15194), .Y(n15192) );
  XNOR2X1 U14713 ( .A(n15195), .B(n15194), .Y(N1576) );
  OAI21X1 U14714 ( .A(n15196), .B(n12827), .C(n15197), .Y(n15194) );
  OAI21X1 U14715 ( .A(N1740), .B(n15198), .C(N1770), .Y(n15197) );
  INVX1 U14716 ( .A(N1740), .Y(n12827) );
  INVX1 U14717 ( .A(n15198), .Y(n15196) );
  XNOR2X1 U14718 ( .A(N1771), .B(N1741), .Y(n15195) );
  XNOR2X1 U14719 ( .A(n15199), .B(n15198), .Y(N1575) );
  OAI21X1 U14720 ( .A(n15200), .B(n12826), .C(n15201), .Y(n15198) );
  OAI21X1 U14721 ( .A(N1739), .B(n15202), .C(N1769), .Y(n15201) );
  INVX1 U14722 ( .A(N1739), .Y(n12826) );
  INVX1 U14723 ( .A(n15202), .Y(n15200) );
  XNOR2X1 U14724 ( .A(N1770), .B(N1740), .Y(n15199) );
  XNOR2X1 U14725 ( .A(n15203), .B(n15202), .Y(N1574) );
  OAI21X1 U14726 ( .A(n15204), .B(n12825), .C(n15205), .Y(n15202) );
  OAI21X1 U14727 ( .A(N1738), .B(n15206), .C(N1768), .Y(n15205) );
  INVX1 U14728 ( .A(N1738), .Y(n12825) );
  INVX1 U14729 ( .A(n15206), .Y(n15204) );
  XNOR2X1 U14730 ( .A(N1769), .B(N1739), .Y(n15203) );
  XNOR2X1 U14731 ( .A(n15207), .B(n15206), .Y(N1573) );
  OAI21X1 U14732 ( .A(n15208), .B(n12824), .C(n15209), .Y(n15206) );
  OAI21X1 U14733 ( .A(N1737), .B(n15210), .C(N1767), .Y(n15209) );
  INVX1 U14734 ( .A(N1737), .Y(n12824) );
  INVX1 U14735 ( .A(n15210), .Y(n15208) );
  XNOR2X1 U14736 ( .A(N1768), .B(N1738), .Y(n15207) );
  XNOR2X1 U14737 ( .A(n15211), .B(n15210), .Y(N1572) );
  OAI21X1 U14738 ( .A(n12823), .B(n15212), .C(n15213), .Y(n15210) );
  OAI21X1 U14739 ( .A(n15214), .B(N1736), .C(N1766), .Y(n15213) );
  INVX1 U14740 ( .A(N1736), .Y(n12823) );
  XNOR2X1 U14741 ( .A(N1767), .B(N1737), .Y(n15211) );
  XNOR2X1 U14742 ( .A(n15214), .B(n15215), .Y(N1571) );
  XNOR2X1 U14743 ( .A(N1766), .B(N1736), .Y(n15215) );
  INVX1 U14744 ( .A(n15212), .Y(n15214) );
  NAND2X1 U14745 ( .A(N1765), .B(N1735), .Y(n15212) );
  XNOR2X1 U14746 ( .A(N1765), .B(n12821), .Y(N1570) );
  INVX1 U14747 ( .A(N1735), .Y(n12821) );
  NOR2X1 U14748 ( .A(n15216), .B(n15217), .Y(N1552) );
  INVX1 U14749 ( .A(N1716), .Y(n15216) );
  XNOR2X1 U14750 ( .A(N1716), .B(n15217), .Y(N1551) );
  NAND2X1 U14751 ( .A(N1715), .B(n15218), .Y(n15217) );
  XOR2X1 U14752 ( .A(n15218), .B(N1715), .Y(N1550) );
  OAI21X1 U14753 ( .A(n15219), .B(n12860), .C(n15220), .Y(n15218) );
  OAI21X1 U14754 ( .A(N1684), .B(n15221), .C(N1714), .Y(n15220) );
  XNOR2X1 U14755 ( .A(n15219), .B(n15222), .Y(N1549) );
  XNOR2X1 U14756 ( .A(N1714), .B(n12860), .Y(n15222) );
  INVX1 U14757 ( .A(N1684), .Y(n12860) );
  INVX1 U14758 ( .A(n15221), .Y(n15219) );
  OAI21X1 U14759 ( .A(n15223), .B(n12859), .C(n15224), .Y(n15221) );
  OAI21X1 U14760 ( .A(N1683), .B(n15225), .C(N1713), .Y(n15224) );
  INVX1 U14761 ( .A(N1683), .Y(n12859) );
  INVX1 U14762 ( .A(n15225), .Y(n15223) );
  XNOR2X1 U14763 ( .A(n15226), .B(n15225), .Y(N1548) );
  OAI21X1 U14764 ( .A(n15227), .B(n12858), .C(n15228), .Y(n15225) );
  OAI21X1 U14765 ( .A(N1682), .B(n15229), .C(N1712), .Y(n15228) );
  INVX1 U14766 ( .A(N1682), .Y(n12858) );
  INVX1 U14767 ( .A(n15229), .Y(n15227) );
  XNOR2X1 U14768 ( .A(N1713), .B(N1683), .Y(n15226) );
  XNOR2X1 U14769 ( .A(n15230), .B(n15229), .Y(N1547) );
  OAI21X1 U14770 ( .A(n15231), .B(n12857), .C(n15232), .Y(n15229) );
  OAI21X1 U14771 ( .A(N1681), .B(n15233), .C(N1711), .Y(n15232) );
  INVX1 U14772 ( .A(N1681), .Y(n12857) );
  INVX1 U14773 ( .A(n15233), .Y(n15231) );
  XNOR2X1 U14774 ( .A(N1712), .B(N1682), .Y(n15230) );
  XNOR2X1 U14775 ( .A(n15234), .B(n15233), .Y(N1546) );
  OAI21X1 U14776 ( .A(n15235), .B(n12856), .C(n15236), .Y(n15233) );
  OAI21X1 U14777 ( .A(N1680), .B(n15237), .C(N1710), .Y(n15236) );
  INVX1 U14778 ( .A(N1680), .Y(n12856) );
  INVX1 U14779 ( .A(n15237), .Y(n15235) );
  XNOR2X1 U14780 ( .A(N1711), .B(N1681), .Y(n15234) );
  XNOR2X1 U14781 ( .A(n15238), .B(n15237), .Y(N1545) );
  OAI21X1 U14782 ( .A(n15239), .B(n12855), .C(n15240), .Y(n15237) );
  OAI21X1 U14783 ( .A(N1679), .B(n15241), .C(N1709), .Y(n15240) );
  INVX1 U14784 ( .A(N1679), .Y(n12855) );
  INVX1 U14785 ( .A(n15241), .Y(n15239) );
  XNOR2X1 U14786 ( .A(N1710), .B(N1680), .Y(n15238) );
  XNOR2X1 U14787 ( .A(n15242), .B(n15241), .Y(N1544) );
  OAI21X1 U14788 ( .A(n12854), .B(n15243), .C(n15244), .Y(n15241) );
  OAI21X1 U14789 ( .A(n15245), .B(N1678), .C(N1708), .Y(n15244) );
  INVX1 U14790 ( .A(N1678), .Y(n12854) );
  XNOR2X1 U14791 ( .A(N1709), .B(N1679), .Y(n15242) );
  XNOR2X1 U14792 ( .A(n15245), .B(n15246), .Y(N1543) );
  XNOR2X1 U14793 ( .A(N1708), .B(N1678), .Y(n15246) );
  INVX1 U14794 ( .A(n15243), .Y(n15245) );
  NAND2X1 U14795 ( .A(N1707), .B(N1677), .Y(n15243) );
  XNOR2X1 U14796 ( .A(N1707), .B(n12852), .Y(N1542) );
  INVX1 U14797 ( .A(N1677), .Y(n12852) );
  NOR2X1 U14798 ( .A(n15247), .B(n15248), .Y(N1522) );
  INVX1 U14799 ( .A(N1656), .Y(n15247) );
  XNOR2X1 U14800 ( .A(N1656), .B(n15248), .Y(N1521) );
  NAND2X1 U14801 ( .A(N1655), .B(n15249), .Y(n15248) );
  XOR2X1 U14802 ( .A(N1655), .B(n15249), .Y(N1520) );
  NOR2X1 U14803 ( .A(n15250), .B(n15251), .Y(n15249) );
  INVX1 U14804 ( .A(N1654), .Y(n15250) );
  XNOR2X1 U14805 ( .A(N1654), .B(n15251), .Y(N1519) );
  NAND2X1 U14806 ( .A(N1653), .B(n15252), .Y(n15251) );
  XOR2X1 U14807 ( .A(n15252), .B(N1653), .Y(N1518) );
  OAI21X1 U14808 ( .A(n15253), .B(n12889), .C(n15254), .Y(n15252) );
  OAI21X1 U14809 ( .A(N1622), .B(n15255), .C(N1652), .Y(n15254) );
  XNOR2X1 U14810 ( .A(n15253), .B(n15256), .Y(N1517) );
  XNOR2X1 U14811 ( .A(N1652), .B(n12889), .Y(n15256) );
  INVX1 U14812 ( .A(N1622), .Y(n12889) );
  INVX1 U14813 ( .A(n15255), .Y(n15253) );
  OAI21X1 U14814 ( .A(n15257), .B(n12888), .C(n15258), .Y(n15255) );
  OAI21X1 U14815 ( .A(N1621), .B(n15259), .C(N1651), .Y(n15258) );
  XNOR2X1 U14816 ( .A(n15257), .B(n15260), .Y(N1516) );
  XNOR2X1 U14817 ( .A(N1651), .B(n12888), .Y(n15260) );
  INVX1 U14818 ( .A(N1621), .Y(n12888) );
  INVX1 U14819 ( .A(n15259), .Y(n15257) );
  OAI21X1 U14820 ( .A(n15261), .B(n12887), .C(n15262), .Y(n15259) );
  OAI21X1 U14821 ( .A(N1620), .B(n15263), .C(N1650), .Y(n15262) );
  INVX1 U14822 ( .A(N1620), .Y(n12887) );
  INVX1 U14823 ( .A(n15263), .Y(n15261) );
  XNOR2X1 U14824 ( .A(n15264), .B(n15263), .Y(N1515) );
  OAI21X1 U14825 ( .A(n15265), .B(n12886), .C(n15266), .Y(n15263) );
  OAI21X1 U14826 ( .A(N1619), .B(n15267), .C(N1649), .Y(n15266) );
  INVX1 U14827 ( .A(N1619), .Y(n12886) );
  INVX1 U14828 ( .A(n15267), .Y(n15265) );
  XNOR2X1 U14829 ( .A(N1650), .B(N1620), .Y(n15264) );
  XNOR2X1 U14830 ( .A(n15268), .B(n15267), .Y(N1514) );
  OAI21X1 U14831 ( .A(n15269), .B(n12885), .C(n15270), .Y(n15267) );
  OAI21X1 U14832 ( .A(N1618), .B(n15271), .C(N1648), .Y(n15270) );
  INVX1 U14833 ( .A(N1618), .Y(n12885) );
  INVX1 U14834 ( .A(n15271), .Y(n15269) );
  XNOR2X1 U14835 ( .A(N1649), .B(N1619), .Y(n15268) );
  XNOR2X1 U14836 ( .A(n15272), .B(n15271), .Y(N1513) );
  OAI21X1 U14837 ( .A(n15273), .B(n12884), .C(n15274), .Y(n15271) );
  OAI21X1 U14838 ( .A(N1617), .B(n15275), .C(N1647), .Y(n15274) );
  INVX1 U14839 ( .A(N1617), .Y(n12884) );
  INVX1 U14840 ( .A(n15275), .Y(n15273) );
  XNOR2X1 U14841 ( .A(N1648), .B(N1618), .Y(n15272) );
  XNOR2X1 U14842 ( .A(n15276), .B(n15275), .Y(N1512) );
  OAI21X1 U14843 ( .A(n12883), .B(n15277), .C(n15278), .Y(n15275) );
  OAI21X1 U14844 ( .A(n15279), .B(N1616), .C(N1646), .Y(n15278) );
  INVX1 U14845 ( .A(N1616), .Y(n12883) );
  XNOR2X1 U14846 ( .A(N1647), .B(N1617), .Y(n15276) );
  XNOR2X1 U14847 ( .A(n15279), .B(n15280), .Y(N1511) );
  XNOR2X1 U14848 ( .A(N1646), .B(N1616), .Y(n15280) );
  INVX1 U14849 ( .A(n15277), .Y(n15279) );
  NAND2X1 U14850 ( .A(N1645), .B(N1615), .Y(n15277) );
  XNOR2X1 U14851 ( .A(N1645), .B(n12881), .Y(N1510) );
  INVX1 U14852 ( .A(N1615), .Y(n12881) );
  XOR2X1 U14853 ( .A(N1417), .B(n15281), .Y(N1402) );
  AND2X1 U14854 ( .A(n15282), .B(N1416), .Y(n15281) );
  XOR2X1 U14855 ( .A(N1416), .B(n15282), .Y(N1401) );
  NOR2X1 U14856 ( .A(n15283), .B(n15284), .Y(n15282) );
  INVX1 U14857 ( .A(N1415), .Y(n15283) );
  XNOR2X1 U14858 ( .A(N1415), .B(n15284), .Y(N1400) );
  NAND2X1 U14859 ( .A(N1414), .B(n15285), .Y(n15284) );
  XOR2X1 U14860 ( .A(N1414), .B(n15285), .Y(N1399) );
  AND2X1 U14861 ( .A(N1413), .B(n15286), .Y(n15285) );
  XOR2X1 U14862 ( .A(n15286), .B(N1413), .Y(N1398) );
  OAI21X1 U14863 ( .A(n15287), .B(n12709), .C(n15288), .Y(n15286) );
  OAI21X1 U14864 ( .A(N1382), .B(n15289), .C(N1412), .Y(n15288) );
  XNOR2X1 U14865 ( .A(n15287), .B(n15290), .Y(N1397) );
  XNOR2X1 U14866 ( .A(N1412), .B(n12709), .Y(n15290) );
  INVX1 U14867 ( .A(N1382), .Y(n12709) );
  INVX1 U14868 ( .A(n15289), .Y(n15287) );
  OAI21X1 U14869 ( .A(n15291), .B(n12708), .C(n15292), .Y(n15289) );
  OAI21X1 U14870 ( .A(N1381), .B(n15293), .C(N1411), .Y(n15292) );
  XNOR2X1 U14871 ( .A(n15291), .B(n15294), .Y(N1396) );
  XNOR2X1 U14872 ( .A(N1411), .B(n12708), .Y(n15294) );
  INVX1 U14873 ( .A(N1381), .Y(n12708) );
  INVX1 U14874 ( .A(n15293), .Y(n15291) );
  OAI21X1 U14875 ( .A(n15295), .B(n12707), .C(n15296), .Y(n15293) );
  OAI21X1 U14876 ( .A(N1380), .B(n15297), .C(N1410), .Y(n15296) );
  INVX1 U14877 ( .A(N1380), .Y(n12707) );
  INVX1 U14878 ( .A(n15297), .Y(n15295) );
  XNOR2X1 U14879 ( .A(n15298), .B(n15297), .Y(N1395) );
  OAI21X1 U14880 ( .A(n15299), .B(n12706), .C(n15300), .Y(n15297) );
  OAI21X1 U14881 ( .A(N1379), .B(n15301), .C(N1409), .Y(n15300) );
  INVX1 U14882 ( .A(N1379), .Y(n12706) );
  INVX1 U14883 ( .A(n15301), .Y(n15299) );
  XNOR2X1 U14884 ( .A(N1410), .B(N1380), .Y(n15298) );
  XNOR2X1 U14885 ( .A(n15302), .B(n15301), .Y(N1394) );
  OAI21X1 U14886 ( .A(n15303), .B(n12705), .C(n15304), .Y(n15301) );
  OAI21X1 U14887 ( .A(N1378), .B(n15305), .C(N1408), .Y(n15304) );
  INVX1 U14888 ( .A(N1378), .Y(n12705) );
  INVX1 U14889 ( .A(n15305), .Y(n15303) );
  XNOR2X1 U14890 ( .A(N1409), .B(N1379), .Y(n15302) );
  XNOR2X1 U14891 ( .A(n15306), .B(n15305), .Y(N1393) );
  OAI21X1 U14892 ( .A(n15307), .B(n12704), .C(n15308), .Y(n15305) );
  OAI21X1 U14893 ( .A(N1377), .B(n15309), .C(N3443), .Y(n15308) );
  INVX1 U14894 ( .A(N1377), .Y(n12704) );
  INVX1 U14895 ( .A(n15309), .Y(n15307) );
  XNOR2X1 U14896 ( .A(N1408), .B(N1378), .Y(n15306) );
  XNOR2X1 U14897 ( .A(n15310), .B(n15309), .Y(N1392) );
  OAI21X1 U14898 ( .A(n12703), .B(n15311), .C(n15312), .Y(n15309) );
  OAI21X1 U14899 ( .A(n15313), .B(N1376), .C(N3442), .Y(n15312) );
  INVX1 U14900 ( .A(n15313), .Y(n15311) );
  INVX1 U14901 ( .A(N1376), .Y(n12703) );
  XNOR2X1 U14902 ( .A(N3443), .B(N1377), .Y(n15310) );
  XNOR2X1 U14903 ( .A(n15313), .B(n15314), .Y(N1391) );
  XNOR2X1 U14904 ( .A(N3442), .B(N1376), .Y(n15314) );
  NOR2X1 U14905 ( .A(n12701), .B(n15162), .Y(n15313) );
  INVX1 U14906 ( .A(N1375), .Y(n12701) );
  XNOR2X1 U14907 ( .A(n15162), .B(N1375), .Y(N1390) );
  INVX1 U14908 ( .A(N3441), .Y(n15162) );
endmodule

