


module WRAP_SRAM ( DataBus, AddressBus, ControlBus, InData, OutData, Address, 
        bCE, bWE, Breq, Bgnt, clk, bReset );
  inout [7:0] DataBus;
  inout [31:0] AddressBus;
  output [7:0] InData;
  input [7:0] OutData;
  output [17:0] Address;
  input Bgnt, clk, bReset;
  output bCE, bWE, Breq;
  inout ControlBus;
  wire   IntEnable, n44, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130;
  tri   [7:0] DataBus;
  tri   AddressBus_31;
  tri   AddressBus_30;
  tri   AddressBus_29;
  tri   AddressBus_28;
  tri   [31:0] AddressBus;
  tri   ControlBus;
  tran( AddressBus_31, AddressBus[31]);
  tran( AddressBus_30, AddressBus[30]);
  tran( AddressBus_29, AddressBus[29]);
  tran( AddressBus_28, AddressBus[28]);

  DFFPOSX1 IntEnable_reg ( .D(n81), .CLK(clk), .Q(IntEnable) );
  DFFPOSX1 \InData_reg[7]  ( .D(n53), .CLK(clk), .Q(InData[7]) );
  DFFPOSX1 \InData_reg[6]  ( .D(n54), .CLK(clk), .Q(InData[6]) );
  DFFPOSX1 \InData_reg[5]  ( .D(n55), .CLK(clk), .Q(InData[5]) );
  DFFPOSX1 \InData_reg[4]  ( .D(n56), .CLK(clk), .Q(InData[4]) );
  DFFPOSX1 \InData_reg[3]  ( .D(n57), .CLK(clk), .Q(InData[3]) );
  DFFPOSX1 \InData_reg[2]  ( .D(n58), .CLK(clk), .Q(InData[2]) );
  DFFPOSX1 \InData_reg[1]  ( .D(n59), .CLK(clk), .Q(InData[1]) );
  DFFPOSX1 \InData_reg[0]  ( .D(n60), .CLK(clk), .Q(InData[0]) );
  DFFPOSX1 \Address_reg[17]  ( .D(n61), .CLK(clk), .Q(Address[17]) );
  DFFPOSX1 \Address_reg[16]  ( .D(n62), .CLK(clk), .Q(Address[16]) );
  DFFPOSX1 \Address_reg[15]  ( .D(n63), .CLK(clk), .Q(Address[15]) );
  DFFPOSX1 \Address_reg[14]  ( .D(n64), .CLK(clk), .Q(Address[14]) );
  DFFPOSX1 \Address_reg[13]  ( .D(n65), .CLK(clk), .Q(Address[13]) );
  DFFPOSX1 \Address_reg[12]  ( .D(n66), .CLK(clk), .Q(Address[12]) );
  DFFPOSX1 \Address_reg[11]  ( .D(n67), .CLK(clk), .Q(Address[11]) );
  DFFPOSX1 \Address_reg[10]  ( .D(n68), .CLK(clk), .Q(Address[10]) );
  DFFPOSX1 \Address_reg[9]  ( .D(n69), .CLK(clk), .Q(Address[9]) );
  DFFPOSX1 \Address_reg[8]  ( .D(n70), .CLK(clk), .Q(Address[8]) );
  DFFPOSX1 \Address_reg[7]  ( .D(n71), .CLK(clk), .Q(Address[7]) );
  DFFPOSX1 \Address_reg[6]  ( .D(n72), .CLK(clk), .Q(Address[6]) );
  DFFPOSX1 \Address_reg[5]  ( .D(n73), .CLK(clk), .Q(Address[5]) );
  DFFPOSX1 \Address_reg[4]  ( .D(n74), .CLK(clk), .Q(Address[4]) );
  DFFPOSX1 \Address_reg[3]  ( .D(n75), .CLK(clk), .Q(Address[3]) );
  DFFPOSX1 \Address_reg[2]  ( .D(n76), .CLK(clk), .Q(Address[2]) );
  DFFPOSX1 \Address_reg[1]  ( .D(n77), .CLK(clk), .Q(Address[1]) );
  DFFPOSX1 \Address_reg[0]  ( .D(n78), .CLK(clk), .Q(Address[0]) );
  DFFPOSX1 bCE_reg ( .D(n79), .CLK(clk), .Q(bCE) );
  DFFPOSX1 bWE_reg ( .D(n80), .CLK(clk), .Q(bWE) );
  DFFPOSX1 Breq_reg ( .D(n52), .CLK(clk), .Q(Breq) );
  TBUFX1 \DataBus_tri[0]  ( .A(n130), .EN(n44), .Y(DataBus[0]) );
  TBUFX1 \DataBus_tri[1]  ( .A(n129), .EN(n44), .Y(DataBus[1]) );
  TBUFX1 \DataBus_tri[2]  ( .A(n128), .EN(n44), .Y(DataBus[2]) );
  TBUFX1 \DataBus_tri[3]  ( .A(n127), .EN(n44), .Y(DataBus[3]) );
  TBUFX1 \DataBus_tri[4]  ( .A(n126), .EN(n44), .Y(DataBus[4]) );
  TBUFX1 \DataBus_tri[5]  ( .A(n125), .EN(n44), .Y(DataBus[5]) );
  TBUFX1 \DataBus_tri[6]  ( .A(n124), .EN(n44), .Y(DataBus[6]) );
  TBUFX1 \DataBus_tri[7]  ( .A(n123), .EN(n44), .Y(DataBus[7]) );
  TBUFX1 ControlBus_tri ( .A(1'b1), .EN(IntEnable), .Y(ControlBus) );
  INVX2 U2 ( .A(n118), .Y(n82) );
  INVX1 U3 ( .A(OutData[7]), .Y(n123) );
  INVX1 U4 ( .A(OutData[6]), .Y(n124) );
  INVX1 U5 ( .A(OutData[5]), .Y(n125) );
  INVX1 U6 ( .A(OutData[4]), .Y(n126) );
  INVX1 U7 ( .A(OutData[3]), .Y(n127) );
  INVX1 U8 ( .A(OutData[2]), .Y(n128) );
  INVX1 U9 ( .A(OutData[1]), .Y(n129) );
  INVX1 U10 ( .A(OutData[0]), .Y(n130) );
  AND2X1 U11 ( .A(bReset), .B(n83), .Y(n81) );
  OAI21X1 U12 ( .A(IntEnable), .B(n84), .C(n82), .Y(n83) );
  INVX1 U13 ( .A(Bgnt), .Y(n84) );
  INVX1 U14 ( .A(n86), .Y(n80) );
  MUX2X1 U15 ( .B(AddressBus[18]), .A(bWE), .S(n82), .Y(n86) );
  INVX1 U16 ( .A(n87), .Y(n79) );
  MUX2X1 U17 ( .B(AddressBus[19]), .A(bCE), .S(n82), .Y(n87) );
  INVX1 U18 ( .A(n88), .Y(n78) );
  MUX2X1 U19 ( .B(AddressBus[0]), .A(Address[0]), .S(n82), .Y(n88) );
  INVX1 U20 ( .A(n89), .Y(n77) );
  MUX2X1 U21 ( .B(AddressBus[1]), .A(Address[1]), .S(n82), .Y(n89) );
  INVX1 U22 ( .A(n90), .Y(n76) );
  MUX2X1 U23 ( .B(AddressBus[2]), .A(Address[2]), .S(n85), .Y(n90) );
  INVX1 U24 ( .A(n91), .Y(n75) );
  MUX2X1 U25 ( .B(AddressBus[3]), .A(Address[3]), .S(n85), .Y(n91) );
  INVX1 U26 ( .A(n92), .Y(n74) );
  MUX2X1 U27 ( .B(AddressBus[4]), .A(Address[4]), .S(n85), .Y(n92) );
  INVX1 U28 ( .A(n93), .Y(n73) );
  MUX2X1 U29 ( .B(AddressBus[5]), .A(Address[5]), .S(n85), .Y(n93) );
  INVX1 U30 ( .A(n94), .Y(n72) );
  MUX2X1 U31 ( .B(AddressBus[6]), .A(Address[6]), .S(n85), .Y(n94) );
  INVX1 U32 ( .A(n95), .Y(n71) );
  MUX2X1 U33 ( .B(AddressBus[7]), .A(Address[7]), .S(n85), .Y(n95) );
  INVX1 U34 ( .A(n96), .Y(n70) );
  MUX2X1 U35 ( .B(AddressBus[8]), .A(Address[8]), .S(n85), .Y(n96) );
  INVX1 U36 ( .A(n97), .Y(n69) );
  MUX2X1 U37 ( .B(AddressBus[9]), .A(Address[9]), .S(n85), .Y(n97) );
  INVX1 U38 ( .A(n98), .Y(n68) );
  MUX2X1 U39 ( .B(AddressBus[10]), .A(Address[10]), .S(n85), .Y(n98) );
  INVX1 U40 ( .A(n99), .Y(n67) );
  MUX2X1 U41 ( .B(AddressBus[11]), .A(Address[11]), .S(n85), .Y(n99) );
  INVX1 U42 ( .A(n100), .Y(n66) );
  MUX2X1 U43 ( .B(AddressBus[12]), .A(Address[12]), .S(n85), .Y(n100) );
  INVX1 U44 ( .A(n101), .Y(n65) );
  MUX2X1 U45 ( .B(AddressBus[13]), .A(Address[13]), .S(n85), .Y(n101) );
  INVX1 U46 ( .A(n102), .Y(n64) );
  MUX2X1 U47 ( .B(AddressBus[14]), .A(Address[14]), .S(n85), .Y(n102) );
  INVX1 U48 ( .A(n103), .Y(n63) );
  MUX2X1 U49 ( .B(AddressBus[15]), .A(Address[15]), .S(n85), .Y(n103) );
  INVX1 U50 ( .A(n104), .Y(n62) );
  MUX2X1 U51 ( .B(AddressBus[16]), .A(Address[16]), .S(n85), .Y(n104) );
  INVX1 U52 ( .A(n105), .Y(n61) );
  MUX2X1 U53 ( .B(AddressBus[17]), .A(Address[17]), .S(n85), .Y(n105) );
  INVX1 U54 ( .A(n106), .Y(n60) );
  MUX2X1 U55 ( .B(DataBus[0]), .A(InData[0]), .S(n85), .Y(n106) );
  INVX1 U56 ( .A(n107), .Y(n59) );
  MUX2X1 U57 ( .B(DataBus[1]), .A(InData[1]), .S(n85), .Y(n107) );
  INVX1 U58 ( .A(n108), .Y(n58) );
  MUX2X1 U59 ( .B(DataBus[2]), .A(InData[2]), .S(n85), .Y(n108) );
  INVX1 U60 ( .A(n109), .Y(n57) );
  MUX2X1 U61 ( .B(DataBus[3]), .A(InData[3]), .S(n85), .Y(n109) );
  INVX1 U62 ( .A(n110), .Y(n56) );
  MUX2X1 U63 ( .B(DataBus[4]), .A(InData[4]), .S(n85), .Y(n110) );
  INVX1 U64 ( .A(n111), .Y(n55) );
  MUX2X1 U65 ( .B(DataBus[5]), .A(InData[5]), .S(n85), .Y(n111) );
  INVX1 U66 ( .A(n112), .Y(n54) );
  MUX2X1 U67 ( .B(DataBus[6]), .A(InData[6]), .S(n85), .Y(n112) );
  INVX1 U68 ( .A(n113), .Y(n53) );
  MUX2X1 U69 ( .B(DataBus[7]), .A(InData[7]), .S(n85), .Y(n113) );
  NOR2X1 U70 ( .A(n114), .B(n115), .Y(n52) );
  INVX1 U71 ( .A(bReset), .Y(n115) );
  AOI22X1 U72 ( .A(n116), .B(n117), .C(Breq), .D(n118), .Y(n114) );
  INVX1 U73 ( .A(n85), .Y(n118) );
  NAND2X1 U74 ( .A(IntEnable), .B(n117), .Y(n85) );
  INVX1 U75 ( .A(n119), .Y(n117) );
  NAND3X1 U76 ( .A(AddressBus_28), .B(n120), .C(n121), .Y(n119) );
  NOR2X1 U77 ( .A(AddressBus_31), .B(AddressBus_30), .Y(n121) );
  INVX1 U78 ( .A(AddressBus_29), .Y(n120) );
  NOR2X1 U79 ( .A(IntEnable), .B(Bgnt), .Y(n116) );
  NOR2X1 U80 ( .A(AddressBus[19]), .B(n122), .Y(n44) );
  INVX1 U81 ( .A(AddressBus[18]), .Y(n122) );
endmodule


module Control_Unit ( Load_XMT_DR, Load_XMT_shftreg, start, shift, clear, 
        Load_XMT_datareg, Byte_ready, T_byte, BC_lt_BCmax, Clock, rst_b );
  input Load_XMT_datareg, Byte_ready, T_byte, BC_lt_BCmax, Clock, rst_b;
  output Load_XMT_DR, Load_XMT_shftreg, start, shift, clear;
  wire   N29, N30, N31, N32, N33, N34, N35, N37, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;
  wire   [2:0] state;
  wire   [2:0] next_state;

  DFFSR \state_reg[0]  ( .D(next_state[0]), .CLK(Clock), .R(1'b1), .S(rst_b), 
        .Q(state[0]) );
  LATCH shift_reg ( .CLK(N29), .D(N30), .Q(shift) );
  LATCH clear_reg ( .CLK(N29), .D(N31), .Q(clear) );
  LATCH \next_state_reg[2]  ( .CLK(N29), .D(N34), .Q(next_state[2]) );
  DFFSR \state_reg[2]  ( .D(next_state[2]), .CLK(Clock), .R(rst_b), .S(1'b1), 
        .Q(state[2]) );
  LATCH \next_state_reg[1]  ( .CLK(N29), .D(N33), .Q(next_state[1]) );
  DFFSR \state_reg[1]  ( .D(next_state[1]), .CLK(Clock), .R(rst_b), .S(1'b1), 
        .Q(state[1]) );
  LATCH \next_state_reg[0]  ( .CLK(N29), .D(N32), .Q(next_state[0]) );
  LATCH Load_XMT_DR_reg ( .CLK(N29), .D(N35), .Q(Load_XMT_DR) );
  LATCH Load_XMT_shftreg_reg ( .CLK(N29), .D(n35), .Q(Load_XMT_shftreg) );
  LATCH start_reg ( .CLK(N29), .D(N37), .Q(start) );
  INVX1 U6 ( .A(n20), .Y(n35) );
  NOR2X1 U7 ( .A(n21), .B(n22), .Y(N35) );
  NAND2X1 U8 ( .A(n23), .B(n24), .Y(n22) );
  OR2X1 U9 ( .A(N37), .B(N30), .Y(N34) );
  NOR2X1 U10 ( .A(n25), .B(n26), .Y(N37) );
  INVX1 U11 ( .A(T_byte), .Y(n25) );
  OAI21X1 U12 ( .A(T_byte), .B(n26), .C(n20), .Y(N33) );
  NAND3X1 U13 ( .A(n23), .B(n21), .C(Byte_ready), .Y(n20) );
  INVX1 U14 ( .A(Load_XMT_datareg), .Y(n21) );
  NAND2X1 U15 ( .A(n27), .B(n28), .Y(N32) );
  OAI21X1 U16 ( .A(Load_XMT_datareg), .B(n24), .C(n23), .Y(n28) );
  INVX1 U17 ( .A(n29), .Y(n23) );
  INVX1 U18 ( .A(Byte_ready), .Y(n24) );
  INVX1 U19 ( .A(N31), .Y(n27) );
  NOR2X1 U20 ( .A(n30), .B(BC_lt_BCmax), .Y(N31) );
  NOR2X1 U21 ( .A(n31), .B(n30), .Y(N30) );
  INVX1 U22 ( .A(BC_lt_BCmax), .Y(n31) );
  NAND3X1 U23 ( .A(n26), .B(n30), .C(n29), .Y(N29) );
  NAND3X1 U24 ( .A(n32), .B(n33), .C(state[0]), .Y(n29) );
  NAND3X1 U25 ( .A(n34), .B(n32), .C(state[2]), .Y(n30) );
  INVX1 U26 ( .A(state[1]), .Y(n32) );
  NAND3X1 U27 ( .A(n34), .B(n33), .C(state[1]), .Y(n26) );
  INVX1 U28 ( .A(state[2]), .Y(n33) );
  INVX1 U29 ( .A(state[0]), .Y(n34) );
endmodule


module Datapath_Unit ( Serial_out, BC_lt_BCmax, Data_Bus, Load_XMT_DR, 
        Load_XMT_shftreg, start, shift, clear, Clock, rst_b );
  input [7:0] Data_Bus;
  input Load_XMT_DR, Load_XMT_shftreg, start, shift, clear, Clock, rst_b;
  output Serial_out, BC_lt_BCmax;
  wire   N55, N56, N57, N58, N59, N60, N61, N62, N63, N81, N82, N84, N85, N87,
         N88, N90, N91, N93, N94, N96, N97, N99, N100, N102, N103, N105, N106,
         N108, N109, N111, N112, N114, N115, N117, N118, N120, N121, N123,
         N124, N126, N127, N129, N130, n127, n128, n130, n84, n129, n131, n132,
         n133, n134, n135, n136, n137, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209;
  wire   [3:0] bit_count;
  tri   Serial_out;
  tri   [8:1] XMT_shftreg;
  tri   [7:0] XMT_datareg;

  DFFSR \XMT_datareg_tri_enable_reg[7]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N82) );
  DFFPOSX1 \XMT_datareg_reg[7]  ( .D(n129), .CLK(Clock), .Q(N81) );
  DFFSR \XMT_datareg_tri_enable_reg[6]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N85) );
  DFFPOSX1 \XMT_datareg_reg[6]  ( .D(n131), .CLK(Clock), .Q(N84) );
  DFFSR \XMT_datareg_tri_enable_reg[5]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N88) );
  DFFPOSX1 \XMT_datareg_reg[5]  ( .D(n132), .CLK(Clock), .Q(N87) );
  DFFSR \XMT_datareg_tri_enable_reg[4]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N91) );
  DFFPOSX1 \XMT_datareg_reg[4]  ( .D(n133), .CLK(Clock), .Q(N90) );
  DFFSR \XMT_datareg_tri_enable_reg[3]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N94) );
  DFFPOSX1 \XMT_datareg_reg[3]  ( .D(n134), .CLK(Clock), .Q(N93) );
  DFFSR \XMT_datareg_tri_enable_reg[2]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N97) );
  DFFPOSX1 \XMT_datareg_reg[2]  ( .D(n135), .CLK(Clock), .Q(N96) );
  DFFSR \XMT_datareg_tri_enable_reg[1]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N100) );
  DFFPOSX1 \XMT_datareg_reg[1]  ( .D(n136), .CLK(Clock), .Q(N99) );
  DFFSR \XMT_datareg_tri_enable_reg[0]  ( .D(1'b0), .CLK(Clock), .R(1'b1), .S(
        rst_b), .Q(N103) );
  DFFPOSX1 \XMT_datareg_reg[0]  ( .D(n137), .CLK(Clock), .Q(N102) );
  DFFSR \XMT_shftreg_tri_enable_reg[8]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N106) );
  DFFSR \XMT_shftreg_reg[8]  ( .D(N63), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N105) );
  DFFSR \XMT_shftreg_tri_enable_reg[7]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N109) );
  DFFSR \XMT_shftreg_reg[7]  ( .D(N62), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N108) );
  DFFSR \XMT_shftreg_tri_enable_reg[6]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N112) );
  DFFSR \XMT_shftreg_reg[6]  ( .D(N61), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N111) );
  DFFSR \XMT_shftreg_tri_enable_reg[5]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N115) );
  DFFSR \XMT_shftreg_reg[5]  ( .D(N60), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N114) );
  DFFSR \XMT_shftreg_tri_enable_reg[4]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N118) );
  DFFSR \XMT_shftreg_reg[4]  ( .D(N59), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N117) );
  DFFSR \XMT_shftreg_tri_enable_reg[3]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N121) );
  DFFSR \XMT_shftreg_reg[3]  ( .D(N58), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N120) );
  DFFSR \XMT_shftreg_tri_enable_reg[2]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N124) );
  DFFSR \XMT_shftreg_reg[2]  ( .D(N57), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N123) );
  DFFSR \XMT_shftreg_tri_enable_reg[1]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N127) );
  DFFSR \XMT_shftreg_reg[1]  ( .D(N56), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N126) );
  DFFSR \XMT_shftreg_tri_enable_reg[0]  ( .D(n84), .CLK(Clock), .R(rst_b), .S(
        1'b1), .Q(N130) );
  DFFSR \XMT_shftreg_reg[0]  ( .D(N55), .CLK(Clock), .R(1'b1), .S(rst_b), .Q(
        N129) );
  DFFSR \bit_count_reg[0]  ( .D(n130), .CLK(Clock), .R(rst_b), .S(1'b1), .Q(
        bit_count[0]) );
  DFFSR \bit_count_reg[1]  ( .D(n127), .CLK(Clock), .R(rst_b), .S(1'b1), .Q(
        bit_count[1]) );
  DFFSR \bit_count_reg[2]  ( .D(n209), .CLK(Clock), .R(rst_b), .S(1'b1), .Q(
        bit_count[2]) );
  DFFSR \bit_count_reg[3]  ( .D(n128), .CLK(Clock), .R(rst_b), .S(1'b1), .Q(
        bit_count[3]) );
  TBUFX1 \XMT_shftreg_tri[0]  ( .A(n208), .EN(n207), .Y(Serial_out) );
  TBUFX1 \XMT_shftreg_tri[1]  ( .A(n206), .EN(n205), .Y(XMT_shftreg[1]) );
  TBUFX1 \XMT_shftreg_tri[2]  ( .A(n204), .EN(n203), .Y(XMT_shftreg[2]) );
  TBUFX1 \XMT_shftreg_tri[3]  ( .A(n202), .EN(n201), .Y(XMT_shftreg[3]) );
  TBUFX1 \XMT_shftreg_tri[4]  ( .A(n200), .EN(n199), .Y(XMT_shftreg[4]) );
  TBUFX1 \XMT_shftreg_tri[5]  ( .A(n198), .EN(n197), .Y(XMT_shftreg[5]) );
  TBUFX1 \XMT_shftreg_tri[6]  ( .A(n196), .EN(n195), .Y(XMT_shftreg[6]) );
  TBUFX1 \XMT_shftreg_tri[7]  ( .A(n194), .EN(n193), .Y(XMT_shftreg[7]) );
  TBUFX1 \XMT_shftreg_tri[8]  ( .A(n192), .EN(n191), .Y(XMT_shftreg[8]) );
  TBUFX1 \XMT_datareg_tri[0]  ( .A(n190), .EN(n189), .Y(XMT_datareg[0]) );
  TBUFX1 \XMT_datareg_tri[1]  ( .A(n188), .EN(n187), .Y(XMT_datareg[1]) );
  TBUFX1 \XMT_datareg_tri[2]  ( .A(n186), .EN(n185), .Y(XMT_datareg[2]) );
  TBUFX1 \XMT_datareg_tri[3]  ( .A(n184), .EN(n183), .Y(XMT_datareg[3]) );
  TBUFX1 \XMT_datareg_tri[4]  ( .A(n182), .EN(n181), .Y(XMT_datareg[4]) );
  TBUFX1 \XMT_datareg_tri[5]  ( .A(n180), .EN(n179), .Y(XMT_datareg[5]) );
  TBUFX1 \XMT_datareg_tri[6]  ( .A(n178), .EN(n177), .Y(XMT_datareg[6]) );
  TBUFX1 \XMT_datareg_tri[7]  ( .A(n176), .EN(n175), .Y(XMT_datareg[7]) );
  INVX1 U3 ( .A(N82), .Y(n175) );
  INVX1 U4 ( .A(N81), .Y(n176) );
  INVX1 U5 ( .A(N85), .Y(n177) );
  INVX1 U6 ( .A(N84), .Y(n178) );
  INVX1 U7 ( .A(N88), .Y(n179) );
  INVX1 U8 ( .A(N87), .Y(n180) );
  INVX1 U9 ( .A(N91), .Y(n181) );
  INVX1 U10 ( .A(N90), .Y(n182) );
  INVX1 U11 ( .A(N94), .Y(n183) );
  INVX1 U12 ( .A(N93), .Y(n184) );
  INVX1 U13 ( .A(N97), .Y(n185) );
  INVX1 U14 ( .A(N96), .Y(n186) );
  INVX1 U15 ( .A(N100), .Y(n187) );
  INVX1 U16 ( .A(N99), .Y(n188) );
  INVX1 U17 ( .A(N103), .Y(n189) );
  INVX1 U18 ( .A(N102), .Y(n190) );
  INVX1 U19 ( .A(N106), .Y(n191) );
  INVX1 U20 ( .A(N105), .Y(n192) );
  INVX1 U21 ( .A(N109), .Y(n193) );
  INVX1 U22 ( .A(N108), .Y(n194) );
  INVX1 U23 ( .A(N112), .Y(n195) );
  INVX1 U24 ( .A(N111), .Y(n196) );
  INVX1 U25 ( .A(N115), .Y(n197) );
  INVX1 U26 ( .A(N114), .Y(n198) );
  INVX1 U27 ( .A(N118), .Y(n199) );
  INVX1 U28 ( .A(N117), .Y(n200) );
  INVX1 U29 ( .A(N121), .Y(n201) );
  INVX1 U30 ( .A(N120), .Y(n202) );
  INVX1 U31 ( .A(N124), .Y(n203) );
  INVX1 U32 ( .A(N123), .Y(n204) );
  INVX1 U33 ( .A(N127), .Y(n205) );
  INVX1 U34 ( .A(N126), .Y(n206) );
  INVX1 U35 ( .A(N130), .Y(n207) );
  INVX1 U36 ( .A(N129), .Y(n208) );
  INVX1 U37 ( .A(n85), .Y(n209) );
  MUX2X1 U38 ( .B(n86), .A(n87), .S(bit_count[2]), .Y(n85) );
  OAI22X1 U39 ( .A(n88), .B(n89), .C(n90), .D(n91), .Y(n84) );
  INVX1 U40 ( .A(n92), .Y(n137) );
  MUX2X1 U41 ( .B(XMT_datareg[0]), .A(Data_Bus[0]), .S(Load_XMT_DR), .Y(n92)
         );
  INVX1 U42 ( .A(n93), .Y(n136) );
  MUX2X1 U43 ( .B(XMT_datareg[1]), .A(Data_Bus[1]), .S(Load_XMT_DR), .Y(n93)
         );
  INVX1 U44 ( .A(n94), .Y(n135) );
  MUX2X1 U45 ( .B(XMT_datareg[2]), .A(Data_Bus[2]), .S(Load_XMT_DR), .Y(n94)
         );
  INVX1 U46 ( .A(n95), .Y(n134) );
  MUX2X1 U47 ( .B(XMT_datareg[3]), .A(Data_Bus[3]), .S(Load_XMT_DR), .Y(n95)
         );
  INVX1 U48 ( .A(n96), .Y(n133) );
  MUX2X1 U49 ( .B(XMT_datareg[4]), .A(Data_Bus[4]), .S(Load_XMT_DR), .Y(n96)
         );
  INVX1 U50 ( .A(n138), .Y(n132) );
  MUX2X1 U51 ( .B(XMT_datareg[5]), .A(Data_Bus[5]), .S(Load_XMT_DR), .Y(n138)
         );
  INVX1 U52 ( .A(n139), .Y(n131) );
  MUX2X1 U53 ( .B(XMT_datareg[6]), .A(Data_Bus[6]), .S(Load_XMT_DR), .Y(n139)
         );
  MUX2X1 U54 ( .B(n140), .A(n141), .S(bit_count[0]), .Y(n130) );
  OR2X1 U55 ( .A(clear), .B(shift), .Y(n141) );
  INVX1 U56 ( .A(n142), .Y(n129) );
  MUX2X1 U57 ( .B(XMT_datareg[7]), .A(Data_Bus[7]), .S(Load_XMT_DR), .Y(n142)
         );
  MUX2X1 U58 ( .B(n143), .A(n144), .S(bit_count[3]), .Y(n128) );
  AOI21X1 U59 ( .A(n145), .B(n146), .C(n87), .Y(n144) );
  OAI21X1 U60 ( .A(bit_count[1]), .B(n140), .C(n147), .Y(n87) );
  INVX1 U61 ( .A(bit_count[2]), .Y(n146) );
  NAND2X1 U62 ( .A(n86), .B(bit_count[2]), .Y(n143) );
  INVX1 U63 ( .A(n148), .Y(n86) );
  NAND3X1 U64 ( .A(bit_count[0]), .B(n145), .C(bit_count[1]), .Y(n148) );
  MUX2X1 U65 ( .B(n149), .A(n147), .S(bit_count[1]), .Y(n127) );
  INVX1 U66 ( .A(n150), .Y(n147) );
  OAI22X1 U67 ( .A(shift), .B(clear), .C(bit_count[0]), .D(n140), .Y(n150) );
  INVX1 U68 ( .A(n145), .Y(n140) );
  NAND2X1 U69 ( .A(bit_count[0]), .B(n145), .Y(n149) );
  NOR2X1 U70 ( .A(n88), .B(clear), .Y(n145) );
  OAI21X1 U71 ( .A(n151), .B(n152), .C(n153), .Y(N63) );
  AOI21X1 U72 ( .A(n154), .B(XMT_datareg[7]), .C(n155), .Y(n153) );
  INVX1 U73 ( .A(n156), .Y(n155) );
  OAI21X1 U74 ( .A(n152), .B(n156), .C(n157), .Y(N62) );
  AOI22X1 U75 ( .A(n154), .B(XMT_datareg[6]), .C(XMT_shftreg[7]), .D(n90), .Y(
        n157) );
  INVX1 U76 ( .A(XMT_shftreg[8]), .Y(n152) );
  OAI21X1 U77 ( .A(n158), .B(n156), .C(n159), .Y(N61) );
  AOI22X1 U78 ( .A(n154), .B(XMT_datareg[5]), .C(XMT_shftreg[6]), .D(n90), .Y(
        n159) );
  INVX1 U79 ( .A(XMT_shftreg[7]), .Y(n158) );
  OAI21X1 U80 ( .A(n156), .B(n160), .C(n161), .Y(N60) );
  AOI22X1 U81 ( .A(n154), .B(XMT_datareg[4]), .C(XMT_shftreg[5]), .D(n90), .Y(
        n161) );
  INVX1 U82 ( .A(XMT_shftreg[6]), .Y(n160) );
  OAI21X1 U83 ( .A(n156), .B(n162), .C(n163), .Y(N59) );
  AOI22X1 U84 ( .A(n154), .B(XMT_datareg[3]), .C(XMT_shftreg[4]), .D(n90), .Y(
        n163) );
  INVX1 U85 ( .A(XMT_shftreg[5]), .Y(n162) );
  OAI21X1 U86 ( .A(n156), .B(n164), .C(n165), .Y(N58) );
  AOI22X1 U87 ( .A(n154), .B(XMT_datareg[2]), .C(XMT_shftreg[3]), .D(n90), .Y(
        n165) );
  INVX1 U88 ( .A(XMT_shftreg[4]), .Y(n164) );
  OAI21X1 U89 ( .A(n156), .B(n166), .C(n167), .Y(N57) );
  AOI22X1 U90 ( .A(n154), .B(XMT_datareg[1]), .C(XMT_shftreg[2]), .D(n90), .Y(
        n167) );
  INVX1 U91 ( .A(XMT_shftreg[3]), .Y(n166) );
  OAI21X1 U92 ( .A(n156), .B(n168), .C(n169), .Y(N56) );
  AOI22X1 U93 ( .A(n154), .B(XMT_datareg[0]), .C(XMT_shftreg[1]), .D(n90), .Y(
        n169) );
  INVX1 U94 ( .A(n151), .Y(n90) );
  INVX1 U95 ( .A(XMT_shftreg[2]), .Y(n168) );
  OAI21X1 U96 ( .A(n156), .B(n170), .C(n171), .Y(N55) );
  AOI21X1 U97 ( .A(n172), .B(Serial_out), .C(n154), .Y(n171) );
  INVX1 U98 ( .A(n173), .Y(n154) );
  NAND3X1 U99 ( .A(n88), .B(n91), .C(Load_XMT_shftreg), .Y(n173) );
  NOR2X1 U100 ( .A(start), .B(n151), .Y(n172) );
  NAND2X1 U101 ( .A(n89), .B(n88), .Y(n151) );
  INVX1 U102 ( .A(shift), .Y(n88) );
  INVX1 U103 ( .A(XMT_shftreg[1]), .Y(n170) );
  NAND3X1 U104 ( .A(n89), .B(n91), .C(shift), .Y(n156) );
  INVX1 U105 ( .A(start), .Y(n91) );
  INVX1 U106 ( .A(Load_XMT_shftreg), .Y(n89) );
  OAI21X1 U107 ( .A(bit_count[0]), .B(n174), .C(bit_count[3]), .Y(BC_lt_BCmax)
         );
  OR2X1 U108 ( .A(bit_count[1]), .B(bit_count[2]), .Y(n174) );
endmodule


module UART_XMTR ( Serial_out, Data_Bus, Load_XMT_datareg, Byte_ready, T_byte, 
        Clock, rst_b );
  input [7:0] Data_Bus;
  input Load_XMT_datareg, Byte_ready, T_byte, Clock, rst_b;
  output Serial_out;
  wire   Load_XMT_DR, Load_XMT_shftreg, start, shift, clear, BC_lt_BCmax;
  tri   Serial_out;

  Control_Unit CONTROL_UNIT_INST ( .Load_XMT_DR(Load_XMT_DR), 
        .Load_XMT_shftreg(Load_XMT_shftreg), .start(start), .shift(shift), 
        .clear(clear), .Load_XMT_datareg(Load_XMT_datareg), .Byte_ready(
        Byte_ready), .T_byte(T_byte), .BC_lt_BCmax(BC_lt_BCmax), .Clock(Clock), 
        .rst_b(rst_b) );
  Datapath_Unit DATAPATH_UNIT_INST ( .Serial_out(Serial_out), .BC_lt_BCmax(
        BC_lt_BCmax), .Data_Bus(Data_Bus), .Load_XMT_DR(Load_XMT_DR), 
        .Load_XMT_shftreg(Load_XMT_shftreg), .start(start), .shift(shift), 
        .clear(clear), .Clock(Clock), .rst_b(rst_b) );
endmodule


module WRAP_UART ( DataBus, AddressBus, ControlBus, InData, Load_XMT_datareg, 
        Byte_ready, T_byte, Breq, Bgnt, clk, bReset );
  inout [7:0] DataBus;
  inout [31:0] AddressBus;
  output [7:0] InData;
  input Bgnt, clk, bReset;
  output Load_XMT_datareg, Byte_ready, T_byte, Breq;
  inout ControlBus;
  wire   IntEnable, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60;
  tri   [7:0] DataBus;
  tri   [31:0] AddressBus;
  tri   AddressBus_2;
  tri   AddressBus_1;
  tri   AddressBus_0;
  tri   ControlBus;
  tran( AddressBus_2, AddressBus[2]);
  tran( AddressBus_1, AddressBus[1]);
  tran( AddressBus_0, AddressBus[0]);

  DFFPOSX1 IntEnable_reg ( .D(n37), .CLK(clk), .Q(IntEnable) );
  DFFPOSX1 Load_XMT_datareg_reg ( .D(n26), .CLK(clk), .Q(Load_XMT_datareg) );
  DFFPOSX1 Byte_ready_reg ( .D(n27), .CLK(clk), .Q(Byte_ready) );
  DFFPOSX1 T_byte_reg ( .D(n28), .CLK(clk), .Q(T_byte) );
  DFFPOSX1 \InData_reg[7]  ( .D(n29), .CLK(clk), .Q(InData[7]) );
  DFFPOSX1 \InData_reg[6]  ( .D(n30), .CLK(clk), .Q(InData[6]) );
  DFFPOSX1 \InData_reg[5]  ( .D(n31), .CLK(clk), .Q(InData[5]) );
  DFFPOSX1 \InData_reg[4]  ( .D(n32), .CLK(clk), .Q(InData[4]) );
  DFFPOSX1 \InData_reg[3]  ( .D(n33), .CLK(clk), .Q(InData[3]) );
  DFFPOSX1 \InData_reg[2]  ( .D(n34), .CLK(clk), .Q(InData[2]) );
  DFFPOSX1 \InData_reg[1]  ( .D(n35), .CLK(clk), .Q(InData[1]) );
  DFFPOSX1 \InData_reg[0]  ( .D(n36), .CLK(clk), .Q(InData[0]) );
  DFFPOSX1 Breq_reg ( .D(n25), .CLK(clk), .Q(Breq) );
  TBUFX1 ControlBus_tri ( .A(1'b1), .EN(IntEnable), .Y(ControlBus) );
  NOR2X1 U3 ( .A(n38), .B(n39), .Y(n37) );
  MUX2X1 U4 ( .B(Bgnt), .A(n40), .S(IntEnable), .Y(n39) );
  INVX1 U5 ( .A(bReset), .Y(n38) );
  INVX1 U6 ( .A(n41), .Y(n36) );
  AOI22X1 U7 ( .A(DataBus[0]), .B(n42), .C(InData[0]), .D(n43), .Y(n41) );
  INVX1 U8 ( .A(n44), .Y(n35) );
  AOI22X1 U9 ( .A(DataBus[1]), .B(n42), .C(InData[1]), .D(n43), .Y(n44) );
  INVX1 U10 ( .A(n45), .Y(n34) );
  AOI22X1 U11 ( .A(DataBus[2]), .B(n42), .C(InData[2]), .D(n43), .Y(n45) );
  INVX1 U12 ( .A(n46), .Y(n33) );
  AOI22X1 U13 ( .A(DataBus[3]), .B(n42), .C(InData[3]), .D(n43), .Y(n46) );
  INVX1 U14 ( .A(n47), .Y(n32) );
  AOI22X1 U15 ( .A(DataBus[4]), .B(n42), .C(InData[4]), .D(n43), .Y(n47) );
  INVX1 U16 ( .A(n48), .Y(n31) );
  AOI22X1 U17 ( .A(DataBus[5]), .B(n42), .C(InData[5]), .D(n43), .Y(n48) );
  INVX1 U18 ( .A(n49), .Y(n30) );
  AOI22X1 U19 ( .A(DataBus[6]), .B(n42), .C(InData[6]), .D(n43), .Y(n49) );
  INVX1 U20 ( .A(n50), .Y(n29) );
  AOI22X1 U21 ( .A(DataBus[7]), .B(n42), .C(InData[7]), .D(n43), .Y(n50) );
  INVX1 U22 ( .A(n51), .Y(n28) );
  AOI22X1 U23 ( .A(AddressBus_2), .B(n42), .C(T_byte), .D(n43), .Y(n51) );
  INVX1 U24 ( .A(n52), .Y(n27) );
  AOI22X1 U25 ( .A(AddressBus_1), .B(n42), .C(Byte_ready), .D(n43), .Y(n52) );
  INVX1 U26 ( .A(n53), .Y(n26) );
  AOI22X1 U27 ( .A(AddressBus_0), .B(n42), .C(Load_XMT_datareg), .D(n43), .Y(
        n53) );
  INVX1 U28 ( .A(n54), .Y(n43) );
  AND2X1 U29 ( .A(IntEnable), .B(n54), .Y(n42) );
  NAND2X1 U30 ( .A(IntEnable), .B(n55), .Y(n54) );
  NOR2X1 U31 ( .A(n56), .B(n57), .Y(n25) );
  NAND2X1 U32 ( .A(n40), .B(bReset), .Y(n57) );
  INVX1 U33 ( .A(n55), .Y(n40) );
  NAND3X1 U34 ( .A(AddressBus[29]), .B(n58), .C(n59), .Y(n55) );
  NOR2X1 U35 ( .A(AddressBus[31]), .B(AddressBus[30]), .Y(n59) );
  INVX1 U36 ( .A(AddressBus[28]), .Y(n58) );
  MUX2X1 U37 ( .B(n60), .A(Breq), .S(IntEnable), .Y(n56) );
  INVX1 U38 ( .A(Bgnt), .Y(n60) );
endmodule


module CannyEdge_DW01_addsub_1 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign B_AS[31] = B[31];
  assign B_AS[30] = B[30];
  assign B_AS[29] = B[29];
  assign B_AS[28] = B[28];
  assign B_AS[27] = B[27];
  assign B_AS[26] = B[26];
  assign B_AS[25] = B[25];
  assign B_AS[24] = B[24];
  assign B_AS[23] = B[23];
  assign B_AS[22] = B[22];
  assign B_AS[21] = B[21];
  assign B_AS[20] = B[20];
  assign B_AS[19] = B[19];
  assign B_AS[18] = B[18];
  assign B_AS[17] = B[17];
  assign B_AS[16] = B[16];
  assign B_AS[15] = B[15];
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_addsub_3 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n24,
         n25, n26, n27, n28, n29, n30;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];

  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  OAI21X1 U10 ( .A(n10), .B(n28), .C(n11), .Y(carry[7]) );
  OAI21X1 U11 ( .A(A[6]), .B(n22), .C(B[6]), .Y(n11) );
  AOI21X1 U12 ( .A(n12), .B(A[5]), .C(n23), .Y(n10) );
  OAI21X1 U13 ( .A(A[5]), .B(n12), .C(B[5]), .Y(n13) );
  OAI21X1 U14 ( .A(n14), .B(n29), .C(n15), .Y(n12) );
  OAI21X1 U15 ( .A(A[4]), .B(n24), .C(B[4]), .Y(n15) );
  AOI21X1 U16 ( .A(n16), .B(A[3]), .C(n25), .Y(n14) );
  OAI21X1 U17 ( .A(A[3]), .B(n16), .C(B[3]), .Y(n17) );
  OAI21X1 U18 ( .A(n18), .B(n30), .C(n19), .Y(n16) );
  OAI21X1 U19 ( .A(A[2]), .B(n26), .C(B[2]), .Y(n19) );
  AOI22X1 U20 ( .A(A[1]), .B(B[1]), .C(B[0]), .D(n27), .Y(n18) );
  OAI21X1 U21 ( .A(A[1]), .B(B[1]), .C(A[0]), .Y(n20) );
  INVX2 U1 ( .A(n10), .Y(n22) );
  INVX2 U2 ( .A(n13), .Y(n23) );
  INVX2 U3 ( .A(n14), .Y(n24) );
  INVX2 U4 ( .A(n17), .Y(n25) );
  INVX2 U5 ( .A(n18), .Y(n26) );
  INVX2 U6 ( .A(n20), .Y(n27) );
  INVX2 U7 ( .A(A[6]), .Y(n28) );
  INVX2 U8 ( .A(A[4]), .Y(n29) );
  INVX2 U9 ( .A(A[2]), .Y(n30) );
endmodule


module CannyEdge_DW01_addsub_4 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign B_AS[14] = B[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_0 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[0] = B[0];

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_1 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_2 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[0] = A[0];
  assign SUM[14] = carry[14];

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_4 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_7 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_8 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_9 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;
  assign SUM[14] = carry[14];

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_10 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_11 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_12 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n16), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n9), .B(B[28]), .Y(n1) );
  AND2X2 U2 ( .A(n10), .B(B[26]), .Y(n2) );
  AND2X2 U3 ( .A(n11), .B(B[24]), .Y(n3) );
  AND2X2 U4 ( .A(n12), .B(B[22]), .Y(n4) );
  AND2X2 U5 ( .A(n13), .B(B[20]), .Y(n5) );
  AND2X2 U6 ( .A(n14), .B(B[18]), .Y(n6) );
  AND2X2 U7 ( .A(n15), .B(B[16]), .Y(n7) );
  AND2X2 U8 ( .A(n1), .B(B[29]), .Y(n8) );
  AND2X2 U9 ( .A(n2), .B(B[27]), .Y(n9) );
  AND2X2 U10 ( .A(n3), .B(B[25]), .Y(n10) );
  AND2X2 U11 ( .A(n4), .B(B[23]), .Y(n11) );
  AND2X2 U12 ( .A(n5), .B(B[21]), .Y(n12) );
  AND2X2 U13 ( .A(n6), .B(B[19]), .Y(n13) );
  AND2X2 U14 ( .A(n7), .B(B[17]), .Y(n14) );
  AND2X2 U15 ( .A(carry[15]), .B(B[15]), .Y(n15) );
  AND2X2 U16 ( .A(B[0]), .B(A[0]), .Y(n16) );
  AND2X2 U17 ( .A(n8), .B(B[30]), .Y(n17) );
  XOR2X1 U18 ( .A(B[31]), .B(n17), .Y(SUM[31]) );
  XOR2X1 U19 ( .A(n8), .B(B[30]), .Y(SUM[30]) );
  XOR2X1 U20 ( .A(n1), .B(B[29]), .Y(SUM[29]) );
  XOR2X1 U21 ( .A(n9), .B(B[28]), .Y(SUM[28]) );
  XOR2X1 U22 ( .A(n2), .B(B[27]), .Y(SUM[27]) );
  XOR2X1 U23 ( .A(n10), .B(B[26]), .Y(SUM[26]) );
  XOR2X1 U24 ( .A(n3), .B(B[25]), .Y(SUM[25]) );
  XOR2X1 U25 ( .A(n11), .B(B[24]), .Y(SUM[24]) );
  XOR2X1 U26 ( .A(n4), .B(B[23]), .Y(SUM[23]) );
  XOR2X1 U27 ( .A(n12), .B(B[22]), .Y(SUM[22]) );
  XOR2X1 U28 ( .A(n5), .B(B[21]), .Y(SUM[21]) );
  XOR2X1 U29 ( .A(n13), .B(B[20]), .Y(SUM[20]) );
  XOR2X1 U30 ( .A(n6), .B(B[19]), .Y(SUM[19]) );
  XOR2X1 U31 ( .A(n14), .B(B[18]), .Y(SUM[18]) );
  XOR2X1 U32 ( .A(n7), .B(B[17]), .Y(SUM[17]) );
  XOR2X1 U33 ( .A(n15), .B(B[16]), .Y(SUM[16]) );
  XOR2X1 U34 ( .A(carry[15]), .B(B[15]), .Y(SUM[15]) );
  XOR2X1 U35 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_13 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1;
  wire   [9:1] carry;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B[1]), .B(A[1]), .Y(n1) );
  AND2X2 U2 ( .A(carry[8]), .B(B[8]), .Y(SUM[9]) );
  XOR2X1 U3 ( .A(carry[8]), .B(B[8]), .Y(SUM[8]) );
  XOR2X1 U4 ( .A(B[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_add_14 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n8), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n10), .B(A[28]), .Y(n1) );
  AND2X2 U2 ( .A(n11), .B(A[26]), .Y(n2) );
  AND2X2 U3 ( .A(n12), .B(A[24]), .Y(n3) );
  AND2X2 U4 ( .A(n13), .B(A[22]), .Y(n4) );
  AND2X2 U5 ( .A(n14), .B(A[20]), .Y(n5) );
  AND2X2 U6 ( .A(n15), .B(A[18]), .Y(n6) );
  AND2X2 U7 ( .A(n16), .B(A[16]), .Y(n7) );
  AND2X2 U8 ( .A(B[0]), .B(A[0]), .Y(n8) );
  AND2X2 U9 ( .A(n1), .B(A[29]), .Y(n9) );
  AND2X2 U10 ( .A(n2), .B(A[27]), .Y(n10) );
  AND2X2 U11 ( .A(n3), .B(A[25]), .Y(n11) );
  AND2X2 U12 ( .A(n4), .B(A[23]), .Y(n12) );
  AND2X2 U13 ( .A(n5), .B(A[21]), .Y(n13) );
  AND2X2 U14 ( .A(n6), .B(A[19]), .Y(n14) );
  AND2X2 U15 ( .A(n7), .B(A[17]), .Y(n15) );
  AND2X2 U16 ( .A(carry[15]), .B(A[15]), .Y(n16) );
  AND2X2 U17 ( .A(n9), .B(A[30]), .Y(n17) );
  XOR2X1 U18 ( .A(A[31]), .B(n17), .Y(SUM[31]) );
  XOR2X1 U19 ( .A(n9), .B(A[30]), .Y(SUM[30]) );
  XOR2X1 U20 ( .A(n1), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U21 ( .A(n10), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U22 ( .A(n2), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U23 ( .A(n11), .B(A[26]), .Y(SUM[26]) );
  XOR2X1 U24 ( .A(n3), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U25 ( .A(n12), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U26 ( .A(n4), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U27 ( .A(n13), .B(A[22]), .Y(SUM[22]) );
  XOR2X1 U28 ( .A(n5), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U29 ( .A(n14), .B(A[20]), .Y(SUM[20]) );
  XOR2X1 U30 ( .A(n6), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U31 ( .A(n15), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U32 ( .A(n7), .B(A[17]), .Y(SUM[17]) );
  XOR2X1 U33 ( .A(n16), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U34 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U35 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_15 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_16 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_17 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YS(SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_18 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [14:1] carry;

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U3 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_addsub_5 ( A, B, CI, ADD_SUB, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [15:0] carry;
  wire   [14:0] B_AS;
  assign SUM[0] = A[0];
  assign SUM[14] = carry[14];
  assign B_AS[13] = B[13];
  assign B_AS[12] = B[12];
  assign B_AS[11] = B[11];
  assign B_AS[10] = B[10];
  assign B_AS[9] = B[9];
  assign B_AS[8] = B[8];
  assign B_AS[7] = B[7];
  assign B_AS[6] = B[6];
  assign B_AS[5] = B[5];
  assign B_AS[4] = B[4];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];

  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(n1), .YC(carry[3]), .YS(SUM[2]) );
  AND2X2 U1 ( .A(B_AS[1]), .B(A[1]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[1]), .B(A[1]), .Y(SUM[1]) );
endmodule


module CannyEdge_DW01_addsub_7 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_31 ( .A(A[31]), .B(B_AS[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B_AS[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B_AS[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B_AS[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B_AS[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B_AS[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B_AS[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B_AS[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B_AS[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B_AS[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B_AS[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B_AS[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B_AS[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B_AS[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B_AS[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B_AS[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B_AS[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B_AS[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B_AS[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B_AS[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B_AS[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  XOR2X1 U1 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[31]), .B(carry[0]), .Y(B_AS[31]) );
  XOR2X1 U9 ( .A(B[30]), .B(carry[0]), .Y(B_AS[30]) );
  XOR2X1 U10 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U11 ( .A(B[29]), .B(carry[0]), .Y(B_AS[29]) );
  XOR2X1 U12 ( .A(B[28]), .B(carry[0]), .Y(B_AS[28]) );
  XOR2X1 U13 ( .A(B[27]), .B(carry[0]), .Y(B_AS[27]) );
  XOR2X1 U14 ( .A(B[26]), .B(carry[0]), .Y(B_AS[26]) );
  XOR2X1 U15 ( .A(B[25]), .B(carry[0]), .Y(B_AS[25]) );
  XOR2X1 U16 ( .A(B[24]), .B(carry[0]), .Y(B_AS[24]) );
  XOR2X1 U17 ( .A(B[23]), .B(carry[0]), .Y(B_AS[23]) );
  XOR2X1 U18 ( .A(B[22]), .B(carry[0]), .Y(B_AS[22]) );
  XOR2X1 U19 ( .A(B[21]), .B(carry[0]), .Y(B_AS[21]) );
  XOR2X1 U20 ( .A(B[20]), .B(carry[0]), .Y(B_AS[20]) );
  XOR2X1 U21 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U22 ( .A(B[19]), .B(carry[0]), .Y(B_AS[19]) );
  XOR2X1 U23 ( .A(B[18]), .B(carry[0]), .Y(B_AS[18]) );
  XOR2X1 U24 ( .A(B[17]), .B(carry[0]), .Y(B_AS[17]) );
  XOR2X1 U25 ( .A(B[16]), .B(carry[0]), .Y(B_AS[16]) );
  XOR2X1 U26 ( .A(B[15]), .B(carry[0]), .Y(B_AS[15]) );
  XOR2X1 U27 ( .A(B[14]), .B(carry[0]), .Y(B_AS[14]) );
  XOR2X1 U28 ( .A(B[13]), .B(carry[0]), .Y(B_AS[13]) );
  XOR2X1 U29 ( .A(B[12]), .B(carry[0]), .Y(B_AS[12]) );
  XOR2X1 U30 ( .A(B[11]), .B(carry[0]), .Y(B_AS[11]) );
  XOR2X1 U31 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U32 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_add_19 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_add_20 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [31:1] carry;

  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n9), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n11), .B(B[28]), .Y(n1) );
  AND2X2 U2 ( .A(n12), .B(B[26]), .Y(n2) );
  AND2X2 U3 ( .A(n13), .B(B[24]), .Y(n3) );
  AND2X2 U4 ( .A(n14), .B(B[22]), .Y(n4) );
  AND2X2 U5 ( .A(n15), .B(B[20]), .Y(n5) );
  AND2X2 U6 ( .A(n16), .B(B[18]), .Y(n6) );
  AND2X2 U7 ( .A(n17), .B(B[16]), .Y(n7) );
  AND2X2 U8 ( .A(n22), .B(B[14]), .Y(n8) );
  AND2X2 U9 ( .A(B[0]), .B(A[0]), .Y(n9) );
  AND2X2 U10 ( .A(n1), .B(B[29]), .Y(n10) );
  AND2X2 U11 ( .A(n2), .B(B[27]), .Y(n11) );
  AND2X2 U12 ( .A(n3), .B(B[25]), .Y(n12) );
  AND2X2 U13 ( .A(n4), .B(B[23]), .Y(n13) );
  AND2X2 U14 ( .A(n5), .B(B[21]), .Y(n14) );
  AND2X2 U15 ( .A(n6), .B(B[19]), .Y(n15) );
  AND2X2 U16 ( .A(n7), .B(B[17]), .Y(n16) );
  AND2X2 U17 ( .A(n8), .B(B[15]), .Y(n17) );
  AND2X2 U18 ( .A(carry[9]), .B(B[9]), .Y(n18) );
  AND2X2 U19 ( .A(n18), .B(B[10]), .Y(n19) );
  AND2X2 U20 ( .A(n19), .B(B[11]), .Y(n20) );
  AND2X2 U21 ( .A(n20), .B(B[12]), .Y(n21) );
  AND2X2 U22 ( .A(n21), .B(B[13]), .Y(n22) );
  AND2X2 U23 ( .A(n10), .B(B[30]), .Y(n23) );
  XOR2X1 U24 ( .A(B[31]), .B(n23), .Y(SUM[31]) );
  XOR2X1 U25 ( .A(n10), .B(B[30]), .Y(SUM[30]) );
  XOR2X1 U26 ( .A(n1), .B(B[29]), .Y(SUM[29]) );
  XOR2X1 U27 ( .A(n11), .B(B[28]), .Y(SUM[28]) );
  XOR2X1 U28 ( .A(n2), .B(B[27]), .Y(SUM[27]) );
  XOR2X1 U29 ( .A(n12), .B(B[26]), .Y(SUM[26]) );
  XOR2X1 U30 ( .A(n3), .B(B[25]), .Y(SUM[25]) );
  XOR2X1 U31 ( .A(n13), .B(B[24]), .Y(SUM[24]) );
  XOR2X1 U32 ( .A(n4), .B(B[23]), .Y(SUM[23]) );
  XOR2X1 U33 ( .A(n14), .B(B[22]), .Y(SUM[22]) );
  XOR2X1 U34 ( .A(n5), .B(B[21]), .Y(SUM[21]) );
  XOR2X1 U35 ( .A(n15), .B(B[20]), .Y(SUM[20]) );
  XOR2X1 U36 ( .A(n6), .B(B[19]), .Y(SUM[19]) );
  XOR2X1 U37 ( .A(n16), .B(B[18]), .Y(SUM[18]) );
  XOR2X1 U38 ( .A(n7), .B(B[17]), .Y(SUM[17]) );
  XOR2X1 U39 ( .A(n17), .B(B[16]), .Y(SUM[16]) );
  XOR2X1 U40 ( .A(n8), .B(B[15]), .Y(SUM[15]) );
  XOR2X1 U41 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U42 ( .A(carry[9]), .B(B[9]), .Y(SUM[9]) );
  XOR2X1 U43 ( .A(n18), .B(B[10]), .Y(SUM[10]) );
  XOR2X1 U44 ( .A(n19), .B(B[11]), .Y(SUM[11]) );
  XOR2X1 U45 ( .A(n20), .B(B[12]), .Y(SUM[12]) );
  XOR2X1 U46 ( .A(n21), .B(B[13]), .Y(SUM[13]) );
  XOR2X1 U47 ( .A(n22), .B(B[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_add_21 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [31:1] carry;

  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n17), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(n9), .B(A[29]), .Y(n1) );
  AND2X2 U2 ( .A(n10), .B(A[27]), .Y(n2) );
  AND2X2 U3 ( .A(n11), .B(A[25]), .Y(n3) );
  AND2X2 U4 ( .A(n12), .B(A[23]), .Y(n4) );
  AND2X2 U5 ( .A(n13), .B(A[21]), .Y(n5) );
  AND2X2 U6 ( .A(n14), .B(A[19]), .Y(n6) );
  AND2X2 U7 ( .A(n15), .B(A[17]), .Y(n7) );
  AND2X2 U8 ( .A(n16), .B(A[15]), .Y(n8) );
  AND2X2 U9 ( .A(n2), .B(A[28]), .Y(n9) );
  AND2X2 U10 ( .A(n3), .B(A[26]), .Y(n10) );
  AND2X2 U11 ( .A(n4), .B(A[24]), .Y(n11) );
  AND2X2 U12 ( .A(n5), .B(A[22]), .Y(n12) );
  AND2X2 U13 ( .A(n6), .B(A[20]), .Y(n13) );
  AND2X2 U14 ( .A(n7), .B(A[18]), .Y(n14) );
  AND2X2 U15 ( .A(n8), .B(A[16]), .Y(n15) );
  AND2X2 U16 ( .A(carry[14]), .B(A[14]), .Y(n16) );
  AND2X2 U17 ( .A(B[0]), .B(A[0]), .Y(n17) );
  AND2X2 U18 ( .A(n1), .B(A[30]), .Y(n18) );
  XOR2X1 U19 ( .A(A[31]), .B(n18), .Y(SUM[31]) );
  XOR2X1 U20 ( .A(n1), .B(A[30]), .Y(SUM[30]) );
  XOR2X1 U21 ( .A(n9), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U22 ( .A(n2), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U23 ( .A(n10), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U24 ( .A(n3), .B(A[26]), .Y(SUM[26]) );
  XOR2X1 U25 ( .A(n11), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U26 ( .A(n4), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U27 ( .A(n12), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U28 ( .A(n5), .B(A[22]), .Y(SUM[22]) );
  XOR2X1 U29 ( .A(n13), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U30 ( .A(n6), .B(A[20]), .Y(SUM[20]) );
  XOR2X1 U31 ( .A(n14), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U32 ( .A(n7), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U33 ( .A(n15), .B(A[17]), .Y(SUM[17]) );
  XOR2X1 U34 ( .A(n8), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U35 ( .A(n16), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U36 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
  XOR2X1 U37 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
endmodule


module CannyEdge_DW01_addsub_9 ( A, B, CI, ADD_SUB, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1;
  wire   [7:0] carry;
  wire   [6:0] B_AS;
  assign B_AS[6] = B[6];
  assign B_AS[3] = B[3];
  assign B_AS[2] = B[2];
  assign B_AS[1] = B[1];
  assign B_AS[0] = B[0];

  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[6]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[6]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B_AS[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B_AS[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CannyEdge_DW01_addsub_11 ( A, B, CI, ADD_SUB, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n5, n6, n7, n8, n9, n10, n12, n13, n14, n15;
  wire   [11:0] carry;
  wire   [10:0] B_AS;

  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YS(SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  OAI21X1 U5 ( .A(n12), .B(n15), .C(n5), .Y(carry[3]) );
  OAI21X1 U6 ( .A(A[2]), .B(n6), .C(n7), .Y(n5) );
  XOR2X1 U7 ( .A(B[2]), .B(ADD_SUB), .Y(n7) );
  OAI21X1 U8 ( .A(n8), .B(n14), .C(n9), .Y(n6) );
  OAI21X1 U9 ( .A(A[1]), .B(n13), .C(n10), .Y(n9) );
  XOR2X1 U10 ( .A(B[1]), .B(ADD_SUB), .Y(n10) );
  MUX2X1 U11 ( .B(ADD_SUB), .A(A[0]), .S(B[0]), .Y(n8) );
  XOR2X1 U12 ( .A(B[9]), .B(ADD_SUB), .Y(B_AS[9]) );
  XOR2X1 U13 ( .A(B[8]), .B(ADD_SUB), .Y(B_AS[8]) );
  XOR2X1 U14 ( .A(B[7]), .B(ADD_SUB), .Y(B_AS[7]) );
  XOR2X1 U15 ( .A(B[6]), .B(ADD_SUB), .Y(B_AS[6]) );
  XOR2X1 U16 ( .A(B[5]), .B(ADD_SUB), .Y(B_AS[5]) );
  XOR2X1 U17 ( .A(B[4]), .B(ADD_SUB), .Y(B_AS[4]) );
  XOR2X1 U18 ( .A(B[3]), .B(ADD_SUB), .Y(B_AS[3]) );
  XOR2X1 U19 ( .A(B[10]), .B(ADD_SUB), .Y(B_AS[10]) );
  INVX2 U1 ( .A(n6), .Y(n12) );
  INVX2 U2 ( .A(n8), .Y(n13) );
  INVX2 U3 ( .A(A[1]), .Y(n14) );
  INVX2 U4 ( .A(A[2]), .Y(n15) );
endmodule


module CannyEdge_DW01_addsub_12 ( A, B, CI, ADD_SUB, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI, ADD_SUB;
  output CO;

  wire   [11:0] carry;
  wire   [10:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_10 ( .A(A[10]), .B(B_AS[10]), .C(carry[10]), .YS(SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B_AS[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9])
         );
  FAX1 U1_8 ( .A(A[8]), .B(B_AS[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8])
         );
  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  XOR2X1 U1 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U9 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U10 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U11 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;
  tri   [31:0] A;

  OAI21X1 U59 ( .A(B[31]), .B(n59), .C(n60), .Y(LT_LE) );
  OAI21X1 U60 ( .A(n120), .B(n61), .C(A[31]), .Y(n60) );
  NAND2X1 U61 ( .A(A[30]), .B(n59), .Y(n61) );
  OAI21X1 U62 ( .A(B[31]), .B(n177), .C(n62), .Y(n59) );
  AOI21X1 U63 ( .A(A[29]), .B(n133), .C(n63), .Y(n62) );
  AOI21X1 U64 ( .A(B[29]), .B(n176), .C(n64), .Y(n63) );
  OAI21X1 U65 ( .A(A[28]), .B(n132), .C(n65), .Y(n64) );
  OAI21X1 U66 ( .A(B[28]), .B(n175), .C(n66), .Y(n65) );
  AOI21X1 U67 ( .A(A[27]), .B(n131), .C(n67), .Y(n66) );
  AOI21X1 U68 ( .A(B[27]), .B(n174), .C(n68), .Y(n67) );
  OAI21X1 U69 ( .A(A[26]), .B(n130), .C(n69), .Y(n68) );
  OAI21X1 U70 ( .A(B[26]), .B(n173), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(A[25]), .B(n129), .C(n71), .Y(n70) );
  AOI21X1 U72 ( .A(B[25]), .B(n172), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(A[24]), .B(n128), .C(n73), .Y(n72) );
  OAI21X1 U74 ( .A(B[24]), .B(n171), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(A[23]), .B(n127), .C(n75), .Y(n74) );
  AOI21X1 U76 ( .A(B[23]), .B(n170), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(A[22]), .B(n126), .C(n77), .Y(n76) );
  OAI21X1 U78 ( .A(B[22]), .B(n169), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(A[21]), .B(n125), .C(n79), .Y(n78) );
  AOI21X1 U80 ( .A(B[21]), .B(n168), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(A[20]), .B(n124), .C(n81), .Y(n80) );
  OAI21X1 U82 ( .A(B[20]), .B(n167), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(A[19]), .B(n123), .C(n83), .Y(n82) );
  AOI21X1 U84 ( .A(B[19]), .B(n166), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(A[18]), .B(n122), .C(n85), .Y(n84) );
  OAI21X1 U86 ( .A(B[18]), .B(n165), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(A[17]), .B(n121), .C(n87), .Y(n86) );
  AOI21X1 U88 ( .A(B[17]), .B(n164), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(A[16]), .B(n134), .C(n89), .Y(n88) );
  OAI21X1 U90 ( .A(B[16]), .B(n163), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(A[15]), .B(n135), .C(n91), .Y(n90) );
  AOI21X1 U92 ( .A(B[15]), .B(n162), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(A[14]), .B(n136), .C(n93), .Y(n92) );
  OAI21X1 U94 ( .A(B[14]), .B(n161), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(A[13]), .B(n137), .C(n95), .Y(n94) );
  AOI21X1 U96 ( .A(B[13]), .B(n160), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(A[12]), .B(n138), .C(n97), .Y(n96) );
  OAI21X1 U98 ( .A(B[12]), .B(n159), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(A[11]), .B(n139), .C(n99), .Y(n98) );
  AOI21X1 U100 ( .A(B[11]), .B(n158), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(A[10]), .B(n140), .C(n101), .Y(n100) );
  OAI21X1 U102 ( .A(B[9]), .B(n157), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(A[10]), .B(n140), .C(n103), .Y(n102) );
  AOI21X1 U104 ( .A(B[9]), .B(n157), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(A[8]), .B(n141), .C(n105), .Y(n104) );
  OAI21X1 U106 ( .A(B[8]), .B(n156), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(A[7]), .B(n142), .C(n107), .Y(n106) );
  AOI21X1 U108 ( .A(B[7]), .B(n155), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(A[6]), .B(n143), .C(n109), .Y(n108) );
  OAI21X1 U110 ( .A(B[6]), .B(n154), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(A[5]), .B(n144), .C(n111), .Y(n110) );
  AOI21X1 U112 ( .A(B[5]), .B(n153), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(A[4]), .B(n145), .C(n113), .Y(n112) );
  OAI21X1 U114 ( .A(B[4]), .B(n152), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(A[3]), .B(n146), .C(n115), .Y(n114) );
  AOI21X1 U116 ( .A(B[3]), .B(n151), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(A[2]), .B(n147), .C(n117), .Y(n116) );
  OAI21X1 U118 ( .A(B[2]), .B(n150), .C(n118), .Y(n117) );
  AOI22X1 U119 ( .A(n119), .B(A[0]), .C(A[1]), .D(n148), .Y(n118) );
  AOI21X1 U120 ( .A(B[1]), .B(n149), .C(B[0]), .Y(n119) );
  INVX2 U1 ( .A(B[31]), .Y(n120) );
  INVX2 U2 ( .A(B[17]), .Y(n121) );
  INVX2 U3 ( .A(B[18]), .Y(n122) );
  INVX2 U4 ( .A(B[19]), .Y(n123) );
  INVX2 U5 ( .A(B[20]), .Y(n124) );
  INVX2 U6 ( .A(B[21]), .Y(n125) );
  INVX2 U7 ( .A(B[22]), .Y(n126) );
  INVX2 U8 ( .A(B[23]), .Y(n127) );
  INVX2 U9 ( .A(B[24]), .Y(n128) );
  INVX2 U10 ( .A(B[25]), .Y(n129) );
  INVX2 U11 ( .A(B[26]), .Y(n130) );
  INVX2 U12 ( .A(B[27]), .Y(n131) );
  INVX2 U13 ( .A(B[28]), .Y(n132) );
  INVX2 U14 ( .A(B[29]), .Y(n133) );
  INVX2 U15 ( .A(B[16]), .Y(n134) );
  INVX2 U16 ( .A(B[15]), .Y(n135) );
  INVX2 U17 ( .A(B[14]), .Y(n136) );
  INVX2 U18 ( .A(B[13]), .Y(n137) );
  INVX2 U19 ( .A(B[12]), .Y(n138) );
  INVX2 U20 ( .A(B[11]), .Y(n139) );
  INVX2 U21 ( .A(B[10]), .Y(n140) );
  INVX2 U22 ( .A(B[8]), .Y(n141) );
  INVX2 U23 ( .A(B[7]), .Y(n142) );
  INVX2 U24 ( .A(B[6]), .Y(n143) );
  INVX2 U25 ( .A(B[5]), .Y(n144) );
  INVX2 U26 ( .A(B[4]), .Y(n145) );
  INVX2 U27 ( .A(B[3]), .Y(n146) );
  INVX2 U28 ( .A(B[2]), .Y(n147) );
  INVX2 U29 ( .A(B[1]), .Y(n148) );
  INVX2 U30 ( .A(A[1]), .Y(n149) );
  INVX2 U31 ( .A(A[2]), .Y(n150) );
  INVX2 U32 ( .A(A[3]), .Y(n151) );
  INVX2 U33 ( .A(A[4]), .Y(n152) );
  INVX2 U34 ( .A(A[5]), .Y(n153) );
  INVX2 U35 ( .A(A[6]), .Y(n154) );
  INVX2 U36 ( .A(A[7]), .Y(n155) );
  INVX2 U37 ( .A(A[8]), .Y(n156) );
  INVX2 U38 ( .A(A[9]), .Y(n157) );
  INVX2 U39 ( .A(A[11]), .Y(n158) );
  INVX2 U40 ( .A(A[12]), .Y(n159) );
  INVX2 U41 ( .A(A[13]), .Y(n160) );
  INVX2 U42 ( .A(A[14]), .Y(n161) );
  INVX2 U43 ( .A(A[15]), .Y(n162) );
  INVX2 U44 ( .A(A[16]), .Y(n163) );
  INVX2 U45 ( .A(A[17]), .Y(n164) );
  INVX2 U46 ( .A(A[18]), .Y(n165) );
  INVX2 U47 ( .A(A[19]), .Y(n166) );
  INVX2 U48 ( .A(A[20]), .Y(n167) );
  INVX2 U49 ( .A(A[21]), .Y(n168) );
  INVX2 U50 ( .A(A[22]), .Y(n169) );
  INVX2 U51 ( .A(A[23]), .Y(n170) );
  INVX2 U52 ( .A(A[24]), .Y(n171) );
  INVX2 U53 ( .A(A[25]), .Y(n172) );
  INVX2 U54 ( .A(A[26]), .Y(n173) );
  INVX2 U55 ( .A(A[27]), .Y(n174) );
  INVX2 U56 ( .A(A[28]), .Y(n175) );
  INVX2 U57 ( .A(A[29]), .Y(n176) );
  INVX2 U58 ( .A(A[30]), .Y(n177) );
endmodule


module CannyEdge_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182;
  tri   [31:0] B;

  OAI21X1 U61 ( .A(n124), .B(n61), .C(n62), .Y(LT_LE) );
  OAI21X1 U62 ( .A(n123), .B(n63), .C(n182), .Y(n62) );
  OAI21X1 U64 ( .A(B[30]), .B(n124), .C(n64), .Y(n61) );
  AOI21X1 U65 ( .A(A[29]), .B(n181), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n137), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n180), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n136), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n179), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n135), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n178), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n134), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n177), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n133), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n176), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n132), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n175), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n131), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n174), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n130), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n173), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n129), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n172), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n128), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n171), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n127), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n170), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n126), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n169), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n125), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n168), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n138), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n167), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n139), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n166), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n140), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n165), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n141), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n164), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n142), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n163), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n143), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n162), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n144), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n162), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n144), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n161), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n145), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n160), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n146), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n159), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n147), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n158), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n148), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n149), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n156), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n150), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n155), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n151), .C(n120), .Y(n119) );
  AOI21X1 U121 ( .A(A[1]), .B(n121), .C(n152), .Y(n120) );
  OAI21X1 U122 ( .A(n121), .B(A[1]), .C(n154), .Y(n122) );
  NAND2X1 U123 ( .A(B[0]), .B(n153), .Y(n121) );
  OR2X2 U63 ( .A(A[31]), .B(B[30]), .Y(n63) );
  INVX2 U1 ( .A(n61), .Y(n123) );
  INVX2 U2 ( .A(A[31]), .Y(n124) );
  INVX2 U3 ( .A(A[17]), .Y(n125) );
  INVX2 U4 ( .A(A[18]), .Y(n126) );
  INVX2 U5 ( .A(A[19]), .Y(n127) );
  INVX2 U6 ( .A(A[20]), .Y(n128) );
  INVX2 U7 ( .A(A[21]), .Y(n129) );
  INVX2 U8 ( .A(A[22]), .Y(n130) );
  INVX2 U9 ( .A(A[23]), .Y(n131) );
  INVX2 U10 ( .A(A[24]), .Y(n132) );
  INVX2 U11 ( .A(A[25]), .Y(n133) );
  INVX2 U12 ( .A(A[26]), .Y(n134) );
  INVX2 U13 ( .A(A[27]), .Y(n135) );
  INVX2 U14 ( .A(A[28]), .Y(n136) );
  INVX2 U15 ( .A(A[29]), .Y(n137) );
  INVX2 U16 ( .A(A[16]), .Y(n138) );
  INVX2 U17 ( .A(A[15]), .Y(n139) );
  INVX2 U18 ( .A(A[14]), .Y(n140) );
  INVX2 U19 ( .A(A[13]), .Y(n141) );
  INVX2 U20 ( .A(A[12]), .Y(n142) );
  INVX2 U21 ( .A(A[11]), .Y(n143) );
  INVX2 U22 ( .A(A[9]), .Y(n144) );
  INVX2 U23 ( .A(A[8]), .Y(n145) );
  INVX2 U24 ( .A(A[7]), .Y(n146) );
  INVX2 U25 ( .A(A[6]), .Y(n147) );
  INVX2 U26 ( .A(A[5]), .Y(n148) );
  INVX2 U27 ( .A(A[4]), .Y(n149) );
  INVX2 U28 ( .A(A[3]), .Y(n150) );
  INVX2 U29 ( .A(A[2]), .Y(n151) );
  INVX2 U30 ( .A(n122), .Y(n152) );
  INVX2 U31 ( .A(A[0]), .Y(n153) );
  INVX2 U32 ( .A(B[1]), .Y(n154) );
  INVX2 U33 ( .A(B[2]), .Y(n155) );
  INVX2 U34 ( .A(B[3]), .Y(n156) );
  INVX2 U35 ( .A(B[4]), .Y(n157) );
  INVX2 U36 ( .A(B[5]), .Y(n158) );
  INVX2 U37 ( .A(B[6]), .Y(n159) );
  INVX2 U38 ( .A(B[7]), .Y(n160) );
  INVX2 U39 ( .A(B[8]), .Y(n161) );
  INVX2 U40 ( .A(B[10]), .Y(n162) );
  INVX2 U41 ( .A(B[11]), .Y(n163) );
  INVX2 U42 ( .A(B[12]), .Y(n164) );
  INVX2 U43 ( .A(B[13]), .Y(n165) );
  INVX2 U44 ( .A(B[14]), .Y(n166) );
  INVX2 U45 ( .A(B[15]), .Y(n167) );
  INVX2 U46 ( .A(B[16]), .Y(n168) );
  INVX2 U47 ( .A(B[17]), .Y(n169) );
  INVX2 U48 ( .A(B[18]), .Y(n170) );
  INVX2 U49 ( .A(B[19]), .Y(n171) );
  INVX2 U50 ( .A(B[20]), .Y(n172) );
  INVX2 U51 ( .A(B[21]), .Y(n173) );
  INVX2 U52 ( .A(B[22]), .Y(n174) );
  INVX2 U53 ( .A(B[23]), .Y(n175) );
  INVX2 U54 ( .A(B[24]), .Y(n176) );
  INVX2 U55 ( .A(B[25]), .Y(n177) );
  INVX2 U56 ( .A(B[26]), .Y(n178) );
  INVX2 U57 ( .A(B[27]), .Y(n179) );
  INVX2 U58 ( .A(B[28]), .Y(n180) );
  INVX2 U59 ( .A(B[29]), .Y(n181) );
  INVX2 U60 ( .A(B[31]), .Y(n182) );
endmodule


module CannyEdge_DW01_cmp2_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182;
  tri   [31:0] B;

  OAI21X1 U61 ( .A(n124), .B(n61), .C(n62), .Y(LT_LE) );
  OAI21X1 U62 ( .A(n123), .B(n63), .C(n182), .Y(n62) );
  OAI21X1 U64 ( .A(B[30]), .B(n124), .C(n64), .Y(n61) );
  AOI21X1 U65 ( .A(A[29]), .B(n181), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n137), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n180), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n136), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n179), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n135), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n178), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n134), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n177), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n133), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n176), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n132), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n175), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n131), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n174), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n130), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n173), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n129), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n172), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n128), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n171), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n127), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n170), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n126), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n169), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n125), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n168), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n138), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n167), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n139), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n166), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n140), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n165), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n141), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n164), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n142), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n163), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n143), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n162), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n144), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n162), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n144), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n161), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n145), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n160), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n146), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n159), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n147), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n158), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n148), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n149), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n156), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n150), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n155), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n151), .C(n120), .Y(n119) );
  AOI21X1 U121 ( .A(A[1]), .B(n121), .C(n152), .Y(n120) );
  OAI21X1 U122 ( .A(n121), .B(A[1]), .C(n154), .Y(n122) );
  NAND2X1 U123 ( .A(B[0]), .B(n153), .Y(n121) );
  OR2X2 U63 ( .A(A[31]), .B(B[30]), .Y(n63) );
  INVX2 U1 ( .A(n61), .Y(n123) );
  INVX2 U2 ( .A(A[31]), .Y(n124) );
  INVX2 U3 ( .A(A[17]), .Y(n125) );
  INVX2 U4 ( .A(A[18]), .Y(n126) );
  INVX2 U5 ( .A(A[19]), .Y(n127) );
  INVX2 U6 ( .A(A[20]), .Y(n128) );
  INVX2 U7 ( .A(A[21]), .Y(n129) );
  INVX2 U8 ( .A(A[22]), .Y(n130) );
  INVX2 U9 ( .A(A[23]), .Y(n131) );
  INVX2 U10 ( .A(A[24]), .Y(n132) );
  INVX2 U11 ( .A(A[25]), .Y(n133) );
  INVX2 U12 ( .A(A[26]), .Y(n134) );
  INVX2 U13 ( .A(A[27]), .Y(n135) );
  INVX2 U14 ( .A(A[28]), .Y(n136) );
  INVX2 U15 ( .A(A[29]), .Y(n137) );
  INVX2 U16 ( .A(A[16]), .Y(n138) );
  INVX2 U17 ( .A(A[15]), .Y(n139) );
  INVX2 U18 ( .A(A[14]), .Y(n140) );
  INVX2 U19 ( .A(A[13]), .Y(n141) );
  INVX2 U20 ( .A(A[12]), .Y(n142) );
  INVX2 U21 ( .A(A[11]), .Y(n143) );
  INVX2 U22 ( .A(A[9]), .Y(n144) );
  INVX2 U23 ( .A(A[8]), .Y(n145) );
  INVX2 U24 ( .A(A[7]), .Y(n146) );
  INVX2 U25 ( .A(A[6]), .Y(n147) );
  INVX2 U26 ( .A(A[5]), .Y(n148) );
  INVX2 U27 ( .A(A[4]), .Y(n149) );
  INVX2 U28 ( .A(A[3]), .Y(n150) );
  INVX2 U29 ( .A(A[2]), .Y(n151) );
  INVX2 U30 ( .A(n122), .Y(n152) );
  INVX2 U31 ( .A(A[0]), .Y(n153) );
  INVX2 U32 ( .A(B[1]), .Y(n154) );
  INVX2 U33 ( .A(B[2]), .Y(n155) );
  INVX2 U34 ( .A(B[3]), .Y(n156) );
  INVX2 U35 ( .A(B[4]), .Y(n157) );
  INVX2 U36 ( .A(B[5]), .Y(n158) );
  INVX2 U37 ( .A(B[6]), .Y(n159) );
  INVX2 U38 ( .A(B[7]), .Y(n160) );
  INVX2 U39 ( .A(B[8]), .Y(n161) );
  INVX2 U40 ( .A(B[10]), .Y(n162) );
  INVX2 U41 ( .A(B[11]), .Y(n163) );
  INVX2 U42 ( .A(B[12]), .Y(n164) );
  INVX2 U43 ( .A(B[13]), .Y(n165) );
  INVX2 U44 ( .A(B[14]), .Y(n166) );
  INVX2 U45 ( .A(B[15]), .Y(n167) );
  INVX2 U46 ( .A(B[16]), .Y(n168) );
  INVX2 U47 ( .A(B[17]), .Y(n169) );
  INVX2 U48 ( .A(B[18]), .Y(n170) );
  INVX2 U49 ( .A(B[19]), .Y(n171) );
  INVX2 U50 ( .A(B[20]), .Y(n172) );
  INVX2 U51 ( .A(B[21]), .Y(n173) );
  INVX2 U52 ( .A(B[22]), .Y(n174) );
  INVX2 U53 ( .A(B[23]), .Y(n175) );
  INVX2 U54 ( .A(B[24]), .Y(n176) );
  INVX2 U55 ( .A(B[25]), .Y(n177) );
  INVX2 U56 ( .A(B[26]), .Y(n178) );
  INVX2 U57 ( .A(B[27]), .Y(n179) );
  INVX2 U58 ( .A(B[28]), .Y(n180) );
  INVX2 U59 ( .A(B[29]), .Y(n181) );
  INVX2 U60 ( .A(B[31]), .Y(n182) );
endmodule


module CannyEdge_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n13), .B(\SUMB[5][5] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n53), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n23), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n30), .B(\SUMB[4][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n26), .B(\SUMB[6][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][2] ), .Y(n11) );
  AND2X2 U11 ( .A(n25), .B(\SUMB[6][3] ), .Y(n12) );
  AND2X2 U12 ( .A(n31), .B(\SUMB[4][5] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[7][4] ), .B(n10), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n9), .B(\SUMB[5][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n21), .B(\SUMB[3][1] ), .Y(n27) );
  AND2X2 U27 ( .A(n15), .B(\SUMB[3][2] ), .Y(n28) );
  AND2X2 U28 ( .A(n16), .B(\SUMB[3][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n17), .B(\SUMB[3][4] ), .Y(n30) );
  AND2X2 U30 ( .A(n18), .B(\SUMB[3][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n20), .B(\ab[3][7] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n12), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n11), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n32), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n11), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n12), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n10), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n21), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n27), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n28), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n29), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n30), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n31), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n6), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n7), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n8), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n9), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n13), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n23), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n24), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n25), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n26), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n32), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n14), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n14), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n22), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n23), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n21), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n20), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n18), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n17), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n16), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(n29), .B(\SUMB[5][5] ), .Y(n3) );
  AND2X2 U3 ( .A(n26), .B(\SUMB[7][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n33), .B(\SUMB[5][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n32), .B(\SUMB[5][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n34), .B(\SUMB[3][1] ), .Y(n7) );
  AND2X2 U7 ( .A(n35), .B(\SUMB[3][2] ), .Y(n8) );
  AND2X2 U8 ( .A(n36), .B(\SUMB[3][3] ), .Y(n9) );
  AND2X2 U9 ( .A(n37), .B(\SUMB[3][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n38), .B(\SUMB[3][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n31), .B(\SUMB[6][4] ), .Y(n12) );
  AND2X2 U12 ( .A(n39), .B(\SUMB[3][6] ), .Y(n13) );
  AND2X2 U13 ( .A(n30), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n12), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n21) );
  XNOR2X1 U21 ( .A(n61), .B(n4), .Y(PRODUCT[9]) );
  AND2X2 U22 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[6][2] ), .Y(n24) );
  AND2X2 U24 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n25) );
  AND2X2 U25 ( .A(n5), .B(\SUMB[6][1] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][3] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][4] ), .Y(n28) );
  AND2X2 U28 ( .A(n11), .B(\SUMB[4][5] ), .Y(n29) );
  AND2X2 U29 ( .A(n27), .B(\SUMB[5][3] ), .Y(n30) );
  AND2X2 U30 ( .A(n28), .B(\SUMB[5][4] ), .Y(n31) );
  AND2X2 U31 ( .A(n8), .B(\SUMB[4][2] ), .Y(n32) );
  AND2X2 U32 ( .A(n7), .B(\SUMB[4][1] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n39) );
  AND2X2 U39 ( .A(n13), .B(n25), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n24), .Y(n42) );
  AND2X2 U42 ( .A(n3), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n26), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n24), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n12), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n34), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n35), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n36), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n37), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n38), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n39), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n7), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n8), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n9), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n10), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n11), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n25), .B(n13), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n33), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n32), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n27), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n28), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n29), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n5), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n6), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n30), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n31), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n3), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n4), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n35), .B(\SUMB[6][4] ), .Y(n3) );
  AND2X2 U3 ( .A(n32), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n41), .B(\SUMB[2][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n36), .B(\SUMB[2][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n37), .B(\SUMB[2][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n38), .B(\SUMB[2][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n39), .B(\SUMB[2][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n40), .B(\SUMB[2][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n27), .B(\SUMB[4][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n33), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n11), .B(n44), .Y(n14) );
  AND2X2 U14 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n21) );
  AND2X2 U21 ( .A(n4), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[3][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][5] ), .Y(n27) );
  AND2X2 U27 ( .A(n23), .B(\SUMB[4][1] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][2] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][3] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][4] ), .Y(n31) );
  AND2X2 U31 ( .A(n28), .B(\SUMB[5][1] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][2] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][3] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][4] ), .Y(n35) );
  AND2X2 U35 ( .A(n15), .B(\SUMB[1][2] ), .Y(n36) );
  AND2X2 U36 ( .A(n21), .B(\SUMB[1][3] ), .Y(n37) );
  AND2X2 U37 ( .A(n16), .B(\SUMB[1][4] ), .Y(n38) );
  AND2X2 U38 ( .A(n17), .B(\SUMB[1][5] ), .Y(n39) );
  AND2X2 U39 ( .A(n18), .B(\SUMB[1][6] ), .Y(n40) );
  AND2X2 U40 ( .A(n20), .B(\SUMB[1][1] ), .Y(n41) );
  AND2X2 U41 ( .A(n19), .B(\ab[1][7] ), .Y(n42) );
  XNOR2X1 U42 ( .A(n61), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U43 ( .A(n10), .B(n42), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][3] ), .B(n13), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][2] ), .B(n12), .Y(n46) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n14), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n14), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n20), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n15), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n21), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n16), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n17), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n18), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n19), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n41), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n36), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n37), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n38), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n39), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n40), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n5), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n6), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n7), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n8), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n9), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n42), .B(n10), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n23), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n24), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n25), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n26), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n27), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n28), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n29), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n30), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n31), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n44), .B(n11), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n32), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n33), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n34), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n35), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n46), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n46), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n45), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n45), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n22), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_4 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n12), .B(\SUMB[5][5] ), .Y(n3) );
  AND2X2 U3 ( .A(n22), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n26), .B(\SUMB[4][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n25), .B(\SUMB[6][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n23), .B(\SUMB[6][2] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][3] ), .Y(n11) );
  AND2X2 U11 ( .A(n30), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(\SUMB[7][4] ), .B(n9), .Y(n13) );
  AND2X2 U13 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(n4), .B(\SUMB[7][1] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[5][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][2] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][3] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][4] ), .Y(n25) );
  AND2X2 U25 ( .A(n14), .B(\SUMB[3][1] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n20), .B(\ab[3][7] ), .Y(n31) );
  XNOR2X1 U31 ( .A(n55), .B(n21), .Y(PRODUCT[9]) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n11), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n10), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n31), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n10), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n11), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n9), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n14), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n26), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n27), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n29), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n5), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n6), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n7), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n8), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n22), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n23), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n24), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n25), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n31), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n13), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n13), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n52), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n53), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n54), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n21), .Y(n36) );
  INVX2 U83 ( .A(n40), .Y(n52) );
  INVX2 U84 ( .A(n44), .Y(n53) );
  INVX2 U85 ( .A(n41), .Y(n54) );
  INVX2 U86 ( .A(\A1[7] ), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_6 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n12), .B(\SUMB[5][5] ), .Y(n3) );
  AND2X2 U3 ( .A(n22), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n26), .B(\SUMB[4][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n25), .B(\SUMB[6][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n23), .B(\SUMB[6][2] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][3] ), .Y(n11) );
  AND2X2 U11 ( .A(n30), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(\SUMB[7][4] ), .B(n9), .Y(n13) );
  AND2X2 U13 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n14) );
  AND2X2 U14 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n19) );
  AND2X2 U19 ( .A(n19), .B(\ab[3][6] ), .Y(n20) );
  AND2X2 U20 ( .A(n4), .B(\SUMB[7][1] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[5][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][2] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][3] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][4] ), .Y(n25) );
  AND2X2 U25 ( .A(n14), .B(\SUMB[3][1] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n20), .B(\ab[3][7] ), .Y(n31) );
  XNOR2X1 U31 ( .A(n53), .B(n21), .Y(PRODUCT[9]) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n11), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n10), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n31), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n10), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n11), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n9), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n14), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n15), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n16), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n17), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n18), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n19), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n26), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n27), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n29), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n20), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n5), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n6), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n7), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n8), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n22), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n23), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n24), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n25), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n31), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n13), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n13), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n21), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_8 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n36), .B(\SUMB[6][4] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n33), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n37), .B(\SUMB[2][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[2][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n39), .B(\SUMB[2][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n40), .B(\SUMB[2][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n41), .B(\SUMB[2][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n42), .B(\SUMB[2][6] ), .Y(n11) );
  AND2X2 U11 ( .A(n28), .B(\SUMB[4][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n35), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(n12), .B(n44), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[3][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[4][4] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][1] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][2] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][3] ), .Y(n35) );
  AND2X2 U35 ( .A(n32), .B(\SUMB[5][4] ), .Y(n36) );
  AND2X2 U36 ( .A(n22), .B(\SUMB[1][1] ), .Y(n37) );
  AND2X2 U37 ( .A(n16), .B(\SUMB[1][2] ), .Y(n38) );
  AND2X2 U38 ( .A(n17), .B(\SUMB[1][3] ), .Y(n39) );
  AND2X2 U39 ( .A(n18), .B(\SUMB[1][4] ), .Y(n40) );
  AND2X2 U40 ( .A(n19), .B(\SUMB[1][5] ), .Y(n41) );
  AND2X2 U41 ( .A(n20), .B(\SUMB[1][6] ), .Y(n42) );
  AND2X2 U42 ( .A(n21), .B(\ab[1][7] ), .Y(n43) );
  AND2X2 U43 ( .A(n11), .B(n43), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][3] ), .B(n14), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][2] ), .B(n13), .Y(n46) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n15), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n15), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n22), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n16), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n17), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n18), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n19), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n20), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n21), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n37), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n38), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n39), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n40), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n41), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n42), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n6), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n7), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n8), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n9), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n10), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n43), .B(n11), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n24), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n25), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n26), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n27), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n28), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n29), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n30), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n31), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n32), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n44), .B(n12), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n33), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n34), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n35), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n36), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n46), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n46), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n45), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n45), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n23), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_9 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n16), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n22), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n21), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n20), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n19), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n18), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n17), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n34), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n35), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n37), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n38), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n39), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n33), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n34), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n35), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n36), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n37), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n38), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n39), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n33), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW02_mult_10 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \B[1] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \A1[9] , \A1[8] , \A1[7] , n3, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n52, n53, n54, n55;
  assign PRODUCT[2] = \B[1] ;
  assign \B[1]  = B[1];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  AND2X2 U2 ( .A(n13), .B(\SUMB[5][5] ), .Y(n3) );
  XNOR2X1 U3 ( .A(n53), .B(n22), .Y(PRODUCT[9]) );
  AND2X2 U4 ( .A(n23), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n27), .B(\SUMB[4][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[4][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n30), .B(\SUMB[4][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n26), .B(\SUMB[6][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n24), .B(\SUMB[6][2] ), .Y(n11) );
  AND2X2 U11 ( .A(n25), .B(\SUMB[6][3] ), .Y(n12) );
  AND2X2 U12 ( .A(n31), .B(\SUMB[4][5] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[7][4] ), .B(n10), .Y(n14) );
  AND2X2 U14 ( .A(\ab[3][0] ), .B(\ab[3][2] ), .Y(n15) );
  AND2X2 U15 ( .A(\B[1] ), .B(\ab[3][3] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[3][2] ), .B(\ab[3][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[3][3] ), .B(\ab[3][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[3][4] ), .B(\ab[3][6] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[3][5] ), .B(\ab[3][7] ), .Y(n20) );
  AND2X2 U20 ( .A(n20), .B(\ab[3][6] ), .Y(n21) );
  AND2X2 U21 ( .A(n5), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n6), .B(\SUMB[5][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n7), .B(\SUMB[5][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n8), .B(\SUMB[5][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n9), .B(\SUMB[5][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n15), .B(\SUMB[3][1] ), .Y(n27) );
  AND2X2 U27 ( .A(n16), .B(\SUMB[3][2] ), .Y(n28) );
  AND2X2 U28 ( .A(n17), .B(\SUMB[3][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n18), .B(\SUMB[3][4] ), .Y(n30) );
  AND2X2 U30 ( .A(n19), .B(\SUMB[3][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n21), .B(\ab[3][7] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][3] ), .B(n12), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][2] ), .B(n11), .Y(n34) );
  AND2X2 U34 ( .A(n3), .B(n32), .Y(n35) );
  XOR2X1 U35 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U36 ( .A(\SUMB[7][2] ), .B(n11), .Y(\A1[7] ) );
  XOR2X1 U37 ( .A(\SUMB[7][3] ), .B(n12), .Y(\A1[8] ) );
  XOR2X1 U38 ( .A(\SUMB[7][4] ), .B(n10), .Y(\A1[9] ) );
  XOR2X1 U39 ( .A(\SUMB[3][1] ), .B(n15), .Y(PRODUCT[4]) );
  XOR2X1 U40 ( .A(\SUMB[3][2] ), .B(n16), .Y(\SUMB[4][1] ) );
  XOR2X1 U41 ( .A(\SUMB[3][3] ), .B(n17), .Y(\SUMB[4][2] ) );
  XOR2X1 U42 ( .A(\SUMB[3][4] ), .B(n18), .Y(\SUMB[4][3] ) );
  XOR2X1 U43 ( .A(\SUMB[3][5] ), .B(n19), .Y(\SUMB[4][4] ) );
  XOR2X1 U44 ( .A(\ab[3][6] ), .B(n20), .Y(\SUMB[4][5] ) );
  XOR2X1 U45 ( .A(\SUMB[4][1] ), .B(n27), .Y(PRODUCT[5]) );
  XOR2X1 U46 ( .A(\SUMB[4][2] ), .B(n28), .Y(\SUMB[5][1] ) );
  XOR2X1 U47 ( .A(\SUMB[4][3] ), .B(n29), .Y(\SUMB[5][2] ) );
  XOR2X1 U48 ( .A(\SUMB[4][4] ), .B(n30), .Y(\SUMB[5][3] ) );
  XOR2X1 U49 ( .A(\SUMB[4][5] ), .B(n31), .Y(\SUMB[5][4] ) );
  XOR2X1 U50 ( .A(\ab[3][7] ), .B(n21), .Y(\SUMB[5][5] ) );
  XOR2X1 U51 ( .A(\SUMB[5][1] ), .B(n6), .Y(PRODUCT[6]) );
  XOR2X1 U52 ( .A(\SUMB[5][2] ), .B(n7), .Y(\SUMB[6][1] ) );
  XOR2X1 U53 ( .A(\SUMB[5][3] ), .B(n8), .Y(\SUMB[6][2] ) );
  XOR2X1 U54 ( .A(\SUMB[5][4] ), .B(n9), .Y(\SUMB[6][3] ) );
  XOR2X1 U55 ( .A(\SUMB[5][5] ), .B(n13), .Y(\SUMB[6][4] ) );
  XOR2X1 U56 ( .A(\SUMB[6][1] ), .B(n23), .Y(PRODUCT[7]) );
  XOR2X1 U57 ( .A(\SUMB[6][2] ), .B(n24), .Y(\SUMB[7][1] ) );
  XOR2X1 U58 ( .A(\SUMB[6][3] ), .B(n25), .Y(\SUMB[7][2] ) );
  XOR2X1 U59 ( .A(\SUMB[6][4] ), .B(n26), .Y(\SUMB[7][3] ) );
  XOR2X1 U60 ( .A(n32), .B(n3), .Y(\SUMB[7][4] ) );
  XOR2X1 U61 ( .A(\ab[3][2] ), .B(\ab[3][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U62 ( .A(\ab[3][3] ), .B(\B[1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U63 ( .A(\ab[3][4] ), .B(\ab[3][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U64 ( .A(\ab[3][5] ), .B(\ab[3][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U65 ( .A(\ab[3][6] ), .B(\ab[3][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U66 ( .A(\ab[3][7] ), .B(\ab[3][5] ), .Y(\SUMB[3][5] ) );
  NOR2X1 U67 ( .A(n14), .B(n35), .Y(n40) );
  NAND2X1 U68 ( .A(n14), .B(n35), .Y(n38) );
  NAND2X1 U69 ( .A(n55), .B(n38), .Y(n37) );
  NOR2X1 U70 ( .A(n34), .B(\A1[8] ), .Y(n41) );
  NAND2X1 U71 ( .A(n34), .B(\A1[8] ), .Y(n42) );
  OAI21X1 U72 ( .A(n36), .B(n41), .C(n42), .Y(n47) );
  NOR2X1 U73 ( .A(n33), .B(\A1[9] ), .Y(n44) );
  AND2X1 U74 ( .A(n33), .B(\A1[9] ), .Y(n45) );
  AOI21X1 U75 ( .A(n47), .B(n54), .C(n45), .Y(n39) );
  XOR2X1 U76 ( .A(n37), .B(n39), .Y(PRODUCT[12]) );
  OAI21X1 U77 ( .A(n40), .B(n39), .C(n38), .Y(PRODUCT[13]) );
  NAND2X1 U78 ( .A(n52), .B(n42), .Y(n43) );
  XOR2X1 U79 ( .A(n43), .B(n36), .Y(PRODUCT[10]) );
  NOR2X1 U80 ( .A(n45), .B(n44), .Y(n46) );
  XOR2X1 U81 ( .A(n47), .B(n46), .Y(PRODUCT[11]) );
  NAND2X1 U82 ( .A(\A1[7] ), .B(n22), .Y(n36) );
  INVX2 U83 ( .A(n41), .Y(n52) );
  INVX2 U84 ( .A(\A1[7] ), .Y(n53) );
  INVX2 U85 ( .A(n44), .Y(n54) );
  INVX2 U86 ( .A(n40), .Y(n55) );
endmodule


module CannyEdge_DW02_mult_11 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [7:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , n3, n4, n5, n6, n7, n8, n9, n22, n20, n18, n16, n14,
         n12, n10, \ab[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[30][1] ,
         \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] ,
         \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[30][0] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] ,
         \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][5] , \CARRYB[25][4] ,
         \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] ,
         \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] ,
         \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][6] ,
         \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] ,
         \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] ,
         \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][6] ,
         \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] ,
         \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] ,
         \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \CARRYB[15][6] ,
         \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] ,
         \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][6] ,
         \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] ,
         \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50;

  AND2X2 U2 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n3) );
  AND2X2 U3 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n4) );
  AND2X2 U4 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n5) );
  AND2X2 U5 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n6) );
  AND2X2 U6 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n7) );
  AND2X2 U7 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n8) );
  AND2X2 U8 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n9) );
  XOR2X1 U24 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U25 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U26 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U27 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U28 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U29 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U30 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  NOR2X1 U41 ( .A(n50), .B(n41), .Y(\ab[1][7] ) );
  NOR2X1 U42 ( .A(n49), .B(n41), .Y(\ab[1][6] ) );
  NOR2X1 U43 ( .A(n48), .B(n41), .Y(\ab[1][5] ) );
  NOR2X1 U44 ( .A(n47), .B(n41), .Y(\ab[1][4] ) );
  NOR2X1 U45 ( .A(n46), .B(n41), .Y(\ab[1][3] ) );
  NOR2X1 U46 ( .A(n45), .B(n41), .Y(\ab[1][2] ) );
  NOR2X1 U47 ( .A(n44), .B(n41), .Y(\ab[1][1] ) );
  NOR2X1 U48 ( .A(n43), .B(n41), .Y(\ab[1][0] ) );
  NOR2X1 U49 ( .A(n50), .B(n42), .Y(\ab[0][7] ) );
  NOR2X1 U50 ( .A(n49), .B(n42), .Y(\ab[0][6] ) );
  NOR2X1 U51 ( .A(n48), .B(n42), .Y(\ab[0][5] ) );
  NOR2X1 U52 ( .A(n47), .B(n42), .Y(\ab[0][4] ) );
  NOR2X1 U53 ( .A(n46), .B(n42), .Y(\ab[0][3] ) );
  NOR2X1 U54 ( .A(n45), .B(n42), .Y(\ab[0][2] ) );
  NOR2X1 U55 ( .A(n44), .B(n42), .Y(\ab[0][1] ) );
  NOR2X1 U56 ( .A(n43), .B(n42), .Y(PRODUCT[0]) );
  FAX1 S4_0 ( .A(n34), .B(\CARRYB[30][0] ), .C(\SUMB[30][1] ), .YS(PRODUCT[31]) );
  FAX1 S1_30_0 ( .A(n34), .B(\CARRYB[29][0] ), .C(\SUMB[29][1] ), .YC(
        \CARRYB[30][0] ), .YS(PRODUCT[30]) );
  FAX1 S1_29_0 ( .A(n34), .B(\CARRYB[28][0] ), .C(\SUMB[28][1] ), .YC(
        \CARRYB[29][0] ), .YS(PRODUCT[29]) );
  FAX1 S1_28_0 ( .A(n34), .B(\CARRYB[27][0] ), .C(\SUMB[27][1] ), .YC(
        \CARRYB[28][0] ), .YS(PRODUCT[28]) );
  FAX1 S1_27_0 ( .A(n34), .B(\CARRYB[26][0] ), .C(\SUMB[26][1] ), .YC(
        \CARRYB[27][0] ), .YS(PRODUCT[27]) );
  FAX1 S1_26_0 ( .A(n34), .B(\CARRYB[25][0] ), .C(\SUMB[25][1] ), .YC(
        \CARRYB[26][0] ), .YS(PRODUCT[26]) );
  FAX1 S1_25_0 ( .A(n34), .B(\CARRYB[24][0] ), .C(\SUMB[24][1] ), .YC(
        \CARRYB[25][0] ), .YS(PRODUCT[25]) );
  FAX1 S1_24_0 ( .A(n34), .B(\CARRYB[23][0] ), .C(\SUMB[23][1] ), .YC(
        \CARRYB[24][0] ), .YS(PRODUCT[24]) );
  FAX1 S1_23_0 ( .A(n34), .B(\CARRYB[22][0] ), .C(\SUMB[22][1] ), .YC(
        \CARRYB[23][0] ), .YS(PRODUCT[23]) );
  FAX1 S1_22_0 ( .A(n34), .B(\CARRYB[21][0] ), .C(\SUMB[21][1] ), .YC(
        \CARRYB[22][0] ), .YS(PRODUCT[22]) );
  FAX1 S1_21_0 ( .A(n34), .B(\CARRYB[20][0] ), .C(\SUMB[20][1] ), .YC(
        \CARRYB[21][0] ), .YS(PRODUCT[21]) );
  FAX1 S1_20_0 ( .A(n34), .B(\CARRYB[19][0] ), .C(\SUMB[19][1] ), .YC(
        \CARRYB[20][0] ), .YS(PRODUCT[20]) );
  FAX1 S1_19_0 ( .A(n34), .B(\CARRYB[18][0] ), .C(\SUMB[18][1] ), .YC(
        \CARRYB[19][0] ), .YS(PRODUCT[19]) );
  FAX1 S1_18_0 ( .A(n34), .B(\CARRYB[17][0] ), .C(\SUMB[17][1] ), .YC(
        \CARRYB[18][0] ), .YS(PRODUCT[18]) );
  FAX1 S1_17_0 ( .A(n34), .B(\CARRYB[16][0] ), .C(\SUMB[16][1] ), .YC(
        \CARRYB[17][0] ), .YS(PRODUCT[17]) );
  FAX1 S1_16_0 ( .A(n34), .B(\CARRYB[15][0] ), .C(\SUMB[15][1] ), .YC(
        \CARRYB[16][0] ), .YS(PRODUCT[16]) );
  FAX1 S1_15_0 ( .A(n34), .B(\CARRYB[14][0] ), .C(\SUMB[14][1] ), .YC(
        \CARRYB[15][0] ), .YS(PRODUCT[15]) );
  FAX1 S1_14_0 ( .A(n34), .B(\CARRYB[13][0] ), .C(\SUMB[13][1] ), .YC(
        \CARRYB[14][0] ), .YS(PRODUCT[14]) );
  FAX1 S1_13_0 ( .A(n34), .B(\CARRYB[12][0] ), .C(\SUMB[12][1] ), .YC(
        \CARRYB[13][0] ), .YS(PRODUCT[13]) );
  FAX1 S1_12_0 ( .A(n34), .B(\CARRYB[11][0] ), .C(\SUMB[11][1] ), .YC(
        \CARRYB[12][0] ), .YS(PRODUCT[12]) );
  FAX1 S1_11_0 ( .A(n34), .B(\CARRYB[10][0] ), .C(\SUMB[10][1] ), .YC(
        \CARRYB[11][0] ), .YS(PRODUCT[11]) );
  FAX1 S1_10_0 ( .A(n34), .B(\CARRYB[9][0] ), .C(\SUMB[9][1] ), .YC(
        \CARRYB[10][0] ), .YS(PRODUCT[10]) );
  FAX1 S1_9_0 ( .A(n34), .B(\CARRYB[8][0] ), .C(\SUMB[8][1] ), .YC(
        \CARRYB[9][0] ), .YS(PRODUCT[9]) );
  FAX1 S1_8_0 ( .A(n34), .B(\CARRYB[7][0] ), .C(\SUMB[7][1] ), .YC(
        \CARRYB[8][0] ), .YS(PRODUCT[8]) );
  FAX1 S1_7_0 ( .A(n34), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(PRODUCT[7]) );
  FAX1 S1_6_0 ( .A(n34), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(PRODUCT[6]) );
  FAX1 S1_5_0 ( .A(n34), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(PRODUCT[5]) );
  FAX1 S1_4_0 ( .A(n34), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(PRODUCT[4]) );
  FAX1 S1_3_0 ( .A(n34), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(PRODUCT[3]) );
  FAX1 S1_2_0 ( .A(n34), .B(n9), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), .YS(
        PRODUCT[2]) );
  NAND2X1 U22 ( .A(B[0]), .B(A[9]), .Y(n22) );
  FAX1 S2_30_1 ( .A(n36), .B(\CARRYB[29][1] ), .C(\SUMB[29][2] ), .YS(
        \SUMB[30][1] ) );
  FAX1 S2_29_1 ( .A(n36), .B(\CARRYB[28][1] ), .C(\SUMB[28][2] ), .YC(
        \CARRYB[29][1] ), .YS(\SUMB[29][1] ) );
  FAX1 S2_28_1 ( .A(n36), .B(\CARRYB[27][1] ), .C(\SUMB[27][2] ), .YC(
        \CARRYB[28][1] ), .YS(\SUMB[28][1] ) );
  FAX1 S2_27_1 ( .A(n36), .B(\CARRYB[26][1] ), .C(\SUMB[26][2] ), .YC(
        \CARRYB[27][1] ), .YS(\SUMB[27][1] ) );
  FAX1 S2_26_1 ( .A(n36), .B(\CARRYB[25][1] ), .C(\SUMB[25][2] ), .YC(
        \CARRYB[26][1] ), .YS(\SUMB[26][1] ) );
  FAX1 S2_25_1 ( .A(n36), .B(\CARRYB[24][1] ), .C(\SUMB[24][2] ), .YC(
        \CARRYB[25][1] ), .YS(\SUMB[25][1] ) );
  FAX1 S2_24_1 ( .A(n36), .B(\CARRYB[23][1] ), .C(\SUMB[23][2] ), .YC(
        \CARRYB[24][1] ), .YS(\SUMB[24][1] ) );
  FAX1 S2_23_1 ( .A(n36), .B(\CARRYB[22][1] ), .C(\SUMB[22][2] ), .YC(
        \CARRYB[23][1] ), .YS(\SUMB[23][1] ) );
  FAX1 S2_22_1 ( .A(n36), .B(\CARRYB[21][1] ), .C(\SUMB[21][2] ), .YC(
        \CARRYB[22][1] ), .YS(\SUMB[22][1] ) );
  FAX1 S2_21_1 ( .A(n36), .B(\CARRYB[20][1] ), .C(\SUMB[20][2] ), .YC(
        \CARRYB[21][1] ), .YS(\SUMB[21][1] ) );
  FAX1 S2_20_1 ( .A(n36), .B(\CARRYB[19][1] ), .C(\SUMB[19][2] ), .YC(
        \CARRYB[20][1] ), .YS(\SUMB[20][1] ) );
  FAX1 S2_19_1 ( .A(n36), .B(\CARRYB[18][1] ), .C(\SUMB[18][2] ), .YC(
        \CARRYB[19][1] ), .YS(\SUMB[19][1] ) );
  FAX1 S2_18_1 ( .A(n36), .B(\CARRYB[17][1] ), .C(\SUMB[17][2] ), .YC(
        \CARRYB[18][1] ), .YS(\SUMB[18][1] ) );
  FAX1 S2_17_1 ( .A(n36), .B(\CARRYB[16][1] ), .C(\SUMB[16][2] ), .YC(
        \CARRYB[17][1] ), .YS(\SUMB[17][1] ) );
  FAX1 S2_16_1 ( .A(n36), .B(\CARRYB[15][1] ), .C(\SUMB[15][2] ), .YC(
        \CARRYB[16][1] ), .YS(\SUMB[16][1] ) );
  FAX1 S2_15_1 ( .A(n36), .B(\CARRYB[14][1] ), .C(\SUMB[14][2] ), .YC(
        \CARRYB[15][1] ), .YS(\SUMB[15][1] ) );
  FAX1 S2_14_1 ( .A(n36), .B(\CARRYB[13][1] ), .C(\SUMB[13][2] ), .YC(
        \CARRYB[14][1] ), .YS(\SUMB[14][1] ) );
  FAX1 S2_13_1 ( .A(n36), .B(\CARRYB[12][1] ), .C(\SUMB[12][2] ), .YC(
        \CARRYB[13][1] ), .YS(\SUMB[13][1] ) );
  FAX1 S2_12_1 ( .A(n36), .B(\CARRYB[11][1] ), .C(\SUMB[11][2] ), .YC(
        \CARRYB[12][1] ), .YS(\SUMB[12][1] ) );
  FAX1 S2_11_1 ( .A(n36), .B(\CARRYB[10][1] ), .C(\SUMB[10][2] ), .YC(
        \CARRYB[11][1] ), .YS(\SUMB[11][1] ) );
  FAX1 S2_10_1 ( .A(n36), .B(\CARRYB[9][1] ), .C(\SUMB[9][2] ), .YC(
        \CARRYB[10][1] ), .YS(\SUMB[10][1] ) );
  FAX1 S2_9_1 ( .A(n36), .B(\CARRYB[8][1] ), .C(\SUMB[8][2] ), .YC(
        \CARRYB[9][1] ), .YS(\SUMB[9][1] ) );
  FAX1 S2_8_1 ( .A(n36), .B(\CARRYB[7][1] ), .C(\SUMB[7][2] ), .YC(
        \CARRYB[8][1] ), .YS(\SUMB[8][1] ) );
  FAX1 S2_7_1 ( .A(n36), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S2_6_1 ( .A(n36), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_5_1 ( .A(n36), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_4_1 ( .A(n36), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_3_1 ( .A(n36), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_2_1 ( .A(n36), .B(n8), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), .YS(
        \SUMB[2][1] ) );
  NAND2X1 U18 ( .A(B[1]), .B(A[9]), .Y(n18) );
  FAX1 S2_29_2 ( .A(n38), .B(\CARRYB[28][2] ), .C(\SUMB[28][3] ), .YS(
        \SUMB[29][2] ) );
  FAX1 S2_28_2 ( .A(n38), .B(\CARRYB[27][2] ), .C(\SUMB[27][3] ), .YC(
        \CARRYB[28][2] ), .YS(\SUMB[28][2] ) );
  FAX1 S2_27_2 ( .A(n38), .B(\CARRYB[26][2] ), .C(\SUMB[26][3] ), .YC(
        \CARRYB[27][2] ), .YS(\SUMB[27][2] ) );
  FAX1 S2_26_2 ( .A(n38), .B(\CARRYB[25][2] ), .C(\SUMB[25][3] ), .YC(
        \CARRYB[26][2] ), .YS(\SUMB[26][2] ) );
  FAX1 S2_25_2 ( .A(n38), .B(\CARRYB[24][2] ), .C(\SUMB[24][3] ), .YC(
        \CARRYB[25][2] ), .YS(\SUMB[25][2] ) );
  FAX1 S2_24_2 ( .A(n38), .B(\CARRYB[23][2] ), .C(\SUMB[23][3] ), .YC(
        \CARRYB[24][2] ), .YS(\SUMB[24][2] ) );
  FAX1 S2_23_2 ( .A(n38), .B(\CARRYB[22][2] ), .C(\SUMB[22][3] ), .YC(
        \CARRYB[23][2] ), .YS(\SUMB[23][2] ) );
  FAX1 S2_22_2 ( .A(n38), .B(\CARRYB[21][2] ), .C(\SUMB[21][3] ), .YC(
        \CARRYB[22][2] ), .YS(\SUMB[22][2] ) );
  FAX1 S2_21_2 ( .A(n38), .B(\CARRYB[20][2] ), .C(\SUMB[20][3] ), .YC(
        \CARRYB[21][2] ), .YS(\SUMB[21][2] ) );
  FAX1 S2_20_2 ( .A(n38), .B(\CARRYB[19][2] ), .C(\SUMB[19][3] ), .YC(
        \CARRYB[20][2] ), .YS(\SUMB[20][2] ) );
  FAX1 S2_19_2 ( .A(n38), .B(\CARRYB[18][2] ), .C(\SUMB[18][3] ), .YC(
        \CARRYB[19][2] ), .YS(\SUMB[19][2] ) );
  FAX1 S2_18_2 ( .A(n38), .B(\CARRYB[17][2] ), .C(\SUMB[17][3] ), .YC(
        \CARRYB[18][2] ), .YS(\SUMB[18][2] ) );
  FAX1 S2_17_2 ( .A(n38), .B(\CARRYB[16][2] ), .C(\SUMB[16][3] ), .YC(
        \CARRYB[17][2] ), .YS(\SUMB[17][2] ) );
  FAX1 S2_16_2 ( .A(n38), .B(\CARRYB[15][2] ), .C(\SUMB[15][3] ), .YC(
        \CARRYB[16][2] ), .YS(\SUMB[16][2] ) );
  FAX1 S2_15_2 ( .A(n38), .B(\CARRYB[14][2] ), .C(\SUMB[14][3] ), .YC(
        \CARRYB[15][2] ), .YS(\SUMB[15][2] ) );
  FAX1 S2_14_2 ( .A(n38), .B(\CARRYB[13][2] ), .C(\SUMB[13][3] ), .YC(
        \CARRYB[14][2] ), .YS(\SUMB[14][2] ) );
  FAX1 S2_13_2 ( .A(n38), .B(\CARRYB[12][2] ), .C(\SUMB[12][3] ), .YC(
        \CARRYB[13][2] ), .YS(\SUMB[13][2] ) );
  FAX1 S2_12_2 ( .A(n38), .B(\CARRYB[11][2] ), .C(\SUMB[11][3] ), .YC(
        \CARRYB[12][2] ), .YS(\SUMB[12][2] ) );
  FAX1 S2_11_2 ( .A(n38), .B(\CARRYB[10][2] ), .C(\SUMB[10][3] ), .YC(
        \CARRYB[11][2] ), .YS(\SUMB[11][2] ) );
  FAX1 S2_10_2 ( .A(n38), .B(\CARRYB[9][2] ), .C(\SUMB[9][3] ), .YC(
        \CARRYB[10][2] ), .YS(\SUMB[10][2] ) );
  FAX1 S2_9_2 ( .A(n38), .B(\CARRYB[8][2] ), .C(\SUMB[8][3] ), .YC(
        \CARRYB[9][2] ), .YS(\SUMB[9][2] ) );
  FAX1 S2_8_2 ( .A(n38), .B(\CARRYB[7][2] ), .C(\SUMB[7][3] ), .YC(
        \CARRYB[8][2] ), .YS(\SUMB[8][2] ) );
  FAX1 S2_7_2 ( .A(n38), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(n38), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_5_2 ( .A(n38), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_4_2 ( .A(n38), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_3_2 ( .A(n38), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_2_2 ( .A(n38), .B(n7), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), .YS(
        \SUMB[2][2] ) );
  NAND2X1 U14 ( .A(B[2]), .B(A[9]), .Y(n14) );
  FAX1 S2_28_3 ( .A(n35), .B(\CARRYB[27][3] ), .C(\SUMB[27][4] ), .YS(
        \SUMB[28][3] ) );
  FAX1 S2_27_3 ( .A(n35), .B(\CARRYB[26][3] ), .C(\SUMB[26][4] ), .YC(
        \CARRYB[27][3] ), .YS(\SUMB[27][3] ) );
  FAX1 S2_26_3 ( .A(n35), .B(\CARRYB[25][3] ), .C(\SUMB[25][4] ), .YC(
        \CARRYB[26][3] ), .YS(\SUMB[26][3] ) );
  FAX1 S2_25_3 ( .A(n35), .B(\CARRYB[24][3] ), .C(\SUMB[24][4] ), .YC(
        \CARRYB[25][3] ), .YS(\SUMB[25][3] ) );
  FAX1 S2_24_3 ( .A(n35), .B(\CARRYB[23][3] ), .C(\SUMB[23][4] ), .YC(
        \CARRYB[24][3] ), .YS(\SUMB[24][3] ) );
  FAX1 S2_23_3 ( .A(n35), .B(\CARRYB[22][3] ), .C(\SUMB[22][4] ), .YC(
        \CARRYB[23][3] ), .YS(\SUMB[23][3] ) );
  FAX1 S2_22_3 ( .A(n35), .B(\CARRYB[21][3] ), .C(\SUMB[21][4] ), .YC(
        \CARRYB[22][3] ), .YS(\SUMB[22][3] ) );
  FAX1 S2_21_3 ( .A(n35), .B(\CARRYB[20][3] ), .C(\SUMB[20][4] ), .YC(
        \CARRYB[21][3] ), .YS(\SUMB[21][3] ) );
  FAX1 S2_20_3 ( .A(n35), .B(\CARRYB[19][3] ), .C(\SUMB[19][4] ), .YC(
        \CARRYB[20][3] ), .YS(\SUMB[20][3] ) );
  FAX1 S2_19_3 ( .A(n35), .B(\CARRYB[18][3] ), .C(\SUMB[18][4] ), .YC(
        \CARRYB[19][3] ), .YS(\SUMB[19][3] ) );
  FAX1 S2_18_3 ( .A(n35), .B(\CARRYB[17][3] ), .C(\SUMB[17][4] ), .YC(
        \CARRYB[18][3] ), .YS(\SUMB[18][3] ) );
  FAX1 S2_17_3 ( .A(n35), .B(\CARRYB[16][3] ), .C(\SUMB[16][4] ), .YC(
        \CARRYB[17][3] ), .YS(\SUMB[17][3] ) );
  FAX1 S2_16_3 ( .A(n35), .B(\CARRYB[15][3] ), .C(\SUMB[15][4] ), .YC(
        \CARRYB[16][3] ), .YS(\SUMB[16][3] ) );
  FAX1 S2_15_3 ( .A(n35), .B(\CARRYB[14][3] ), .C(\SUMB[14][4] ), .YC(
        \CARRYB[15][3] ), .YS(\SUMB[15][3] ) );
  FAX1 S2_14_3 ( .A(n35), .B(\CARRYB[13][3] ), .C(\SUMB[13][4] ), .YC(
        \CARRYB[14][3] ), .YS(\SUMB[14][3] ) );
  FAX1 S2_13_3 ( .A(n35), .B(\CARRYB[12][3] ), .C(\SUMB[12][4] ), .YC(
        \CARRYB[13][3] ), .YS(\SUMB[13][3] ) );
  FAX1 S2_12_3 ( .A(n35), .B(\CARRYB[11][3] ), .C(\SUMB[11][4] ), .YC(
        \CARRYB[12][3] ), .YS(\SUMB[12][3] ) );
  FAX1 S2_11_3 ( .A(n35), .B(\CARRYB[10][3] ), .C(\SUMB[10][4] ), .YC(
        \CARRYB[11][3] ), .YS(\SUMB[11][3] ) );
  FAX1 S2_10_3 ( .A(n35), .B(\CARRYB[9][3] ), .C(\SUMB[9][4] ), .YC(
        \CARRYB[10][3] ), .YS(\SUMB[10][3] ) );
  FAX1 S2_9_3 ( .A(n35), .B(\CARRYB[8][3] ), .C(\SUMB[8][4] ), .YC(
        \CARRYB[9][3] ), .YS(\SUMB[9][3] ) );
  FAX1 S2_8_3 ( .A(n35), .B(\CARRYB[7][3] ), .C(\SUMB[7][4] ), .YC(
        \CARRYB[8][3] ), .YS(\SUMB[8][3] ) );
  FAX1 S2_7_3 ( .A(n35), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(n35), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(n35), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_4_3 ( .A(n35), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_3_3 ( .A(n35), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_2_3 ( .A(n35), .B(n6), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), .YS(
        \SUMB[2][3] ) );
  NAND2X1 U20 ( .A(B[3]), .B(A[9]), .Y(n20) );
  FAX1 S2_27_4 ( .A(n37), .B(\CARRYB[26][4] ), .C(\SUMB[26][5] ), .YS(
        \SUMB[27][4] ) );
  FAX1 S2_26_4 ( .A(n37), .B(\CARRYB[25][4] ), .C(\SUMB[25][5] ), .YC(
        \CARRYB[26][4] ), .YS(\SUMB[26][4] ) );
  FAX1 S2_25_4 ( .A(n37), .B(\CARRYB[24][4] ), .C(\SUMB[24][5] ), .YC(
        \CARRYB[25][4] ), .YS(\SUMB[25][4] ) );
  FAX1 S2_24_4 ( .A(n37), .B(\CARRYB[23][4] ), .C(\SUMB[23][5] ), .YC(
        \CARRYB[24][4] ), .YS(\SUMB[24][4] ) );
  FAX1 S2_23_4 ( .A(n37), .B(\CARRYB[22][4] ), .C(\SUMB[22][5] ), .YC(
        \CARRYB[23][4] ), .YS(\SUMB[23][4] ) );
  FAX1 S2_22_4 ( .A(n37), .B(\CARRYB[21][4] ), .C(\SUMB[21][5] ), .YC(
        \CARRYB[22][4] ), .YS(\SUMB[22][4] ) );
  FAX1 S2_21_4 ( .A(n37), .B(\CARRYB[20][4] ), .C(\SUMB[20][5] ), .YC(
        \CARRYB[21][4] ), .YS(\SUMB[21][4] ) );
  FAX1 S2_20_4 ( .A(n37), .B(\CARRYB[19][4] ), .C(\SUMB[19][5] ), .YC(
        \CARRYB[20][4] ), .YS(\SUMB[20][4] ) );
  FAX1 S2_19_4 ( .A(n37), .B(\CARRYB[18][4] ), .C(\SUMB[18][5] ), .YC(
        \CARRYB[19][4] ), .YS(\SUMB[19][4] ) );
  FAX1 S2_18_4 ( .A(n37), .B(\CARRYB[17][4] ), .C(\SUMB[17][5] ), .YC(
        \CARRYB[18][4] ), .YS(\SUMB[18][4] ) );
  FAX1 S2_17_4 ( .A(n37), .B(\CARRYB[16][4] ), .C(\SUMB[16][5] ), .YC(
        \CARRYB[17][4] ), .YS(\SUMB[17][4] ) );
  FAX1 S2_16_4 ( .A(n37), .B(\CARRYB[15][4] ), .C(\SUMB[15][5] ), .YC(
        \CARRYB[16][4] ), .YS(\SUMB[16][4] ) );
  FAX1 S2_15_4 ( .A(n37), .B(\CARRYB[14][4] ), .C(\SUMB[14][5] ), .YC(
        \CARRYB[15][4] ), .YS(\SUMB[15][4] ) );
  FAX1 S2_14_4 ( .A(n37), .B(\CARRYB[13][4] ), .C(\SUMB[13][5] ), .YC(
        \CARRYB[14][4] ), .YS(\SUMB[14][4] ) );
  FAX1 S2_13_4 ( .A(n37), .B(\CARRYB[12][4] ), .C(\SUMB[12][5] ), .YC(
        \CARRYB[13][4] ), .YS(\SUMB[13][4] ) );
  FAX1 S2_12_4 ( .A(n37), .B(\CARRYB[11][4] ), .C(\SUMB[11][5] ), .YC(
        \CARRYB[12][4] ), .YS(\SUMB[12][4] ) );
  FAX1 S2_11_4 ( .A(n37), .B(\CARRYB[10][4] ), .C(\SUMB[10][5] ), .YC(
        \CARRYB[11][4] ), .YS(\SUMB[11][4] ) );
  FAX1 S2_10_4 ( .A(n37), .B(\CARRYB[9][4] ), .C(\SUMB[9][5] ), .YC(
        \CARRYB[10][4] ), .YS(\SUMB[10][4] ) );
  FAX1 S2_9_4 ( .A(n37), .B(\CARRYB[8][4] ), .C(\SUMB[8][5] ), .YC(
        \CARRYB[9][4] ), .YS(\SUMB[9][4] ) );
  FAX1 S2_8_4 ( .A(n37), .B(\CARRYB[7][4] ), .C(\SUMB[7][5] ), .YC(
        \CARRYB[8][4] ), .YS(\SUMB[8][4] ) );
  FAX1 S2_7_4 ( .A(n37), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(n37), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(n37), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(n37), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_3_4 ( .A(n37), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_2_4 ( .A(n37), .B(n5), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), .YS(
        \SUMB[2][4] ) );
  NAND2X1 U16 ( .A(B[4]), .B(A[9]), .Y(n16) );
  FAX1 S2_26_5 ( .A(n39), .B(\CARRYB[25][5] ), .C(\SUMB[25][6] ), .YS(
        \SUMB[26][5] ) );
  FAX1 S3_25_6 ( .A(n40), .B(\CARRYB[24][6] ), .C(\ab[9][7] ), .YS(
        \SUMB[25][6] ) );
  FAX1 S2_25_5 ( .A(n39), .B(\CARRYB[24][5] ), .C(\SUMB[24][6] ), .YC(
        \CARRYB[25][5] ), .YS(\SUMB[25][5] ) );
  FAX1 S3_24_6 ( .A(n40), .B(\CARRYB[23][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[24][6] ), .YS(\SUMB[24][6] ) );
  FAX1 S2_24_5 ( .A(n39), .B(\CARRYB[23][5] ), .C(\SUMB[23][6] ), .YC(
        \CARRYB[24][5] ), .YS(\SUMB[24][5] ) );
  FAX1 S3_23_6 ( .A(n40), .B(\CARRYB[22][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[23][6] ), .YS(\SUMB[23][6] ) );
  FAX1 S2_23_5 ( .A(n39), .B(\CARRYB[22][5] ), .C(\SUMB[22][6] ), .YC(
        \CARRYB[23][5] ), .YS(\SUMB[23][5] ) );
  FAX1 S3_22_6 ( .A(n40), .B(\CARRYB[21][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[22][6] ), .YS(\SUMB[22][6] ) );
  FAX1 S2_22_5 ( .A(n39), .B(\CARRYB[21][5] ), .C(\SUMB[21][6] ), .YC(
        \CARRYB[22][5] ), .YS(\SUMB[22][5] ) );
  FAX1 S3_21_6 ( .A(n40), .B(\CARRYB[20][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[21][6] ), .YS(\SUMB[21][6] ) );
  FAX1 S2_21_5 ( .A(n39), .B(\CARRYB[20][5] ), .C(\SUMB[20][6] ), .YC(
        \CARRYB[21][5] ), .YS(\SUMB[21][5] ) );
  FAX1 S3_20_6 ( .A(n40), .B(\CARRYB[19][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[20][6] ), .YS(\SUMB[20][6] ) );
  FAX1 S2_20_5 ( .A(n39), .B(\CARRYB[19][5] ), .C(\SUMB[19][6] ), .YC(
        \CARRYB[20][5] ), .YS(\SUMB[20][5] ) );
  FAX1 S3_19_6 ( .A(n40), .B(\CARRYB[18][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[19][6] ), .YS(\SUMB[19][6] ) );
  FAX1 S2_19_5 ( .A(n39), .B(\CARRYB[18][5] ), .C(\SUMB[18][6] ), .YC(
        \CARRYB[19][5] ), .YS(\SUMB[19][5] ) );
  FAX1 S3_18_6 ( .A(n40), .B(\CARRYB[17][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[18][6] ), .YS(\SUMB[18][6] ) );
  FAX1 S2_18_5 ( .A(n39), .B(\CARRYB[17][5] ), .C(\SUMB[17][6] ), .YC(
        \CARRYB[18][5] ), .YS(\SUMB[18][5] ) );
  FAX1 S3_17_6 ( .A(n40), .B(\CARRYB[16][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[17][6] ), .YS(\SUMB[17][6] ) );
  FAX1 S2_17_5 ( .A(n39), .B(\CARRYB[16][5] ), .C(\SUMB[16][6] ), .YC(
        \CARRYB[17][5] ), .YS(\SUMB[17][5] ) );
  FAX1 S3_16_6 ( .A(n40), .B(\CARRYB[15][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[16][6] ), .YS(\SUMB[16][6] ) );
  FAX1 S2_16_5 ( .A(n39), .B(\CARRYB[15][5] ), .C(\SUMB[15][6] ), .YC(
        \CARRYB[16][5] ), .YS(\SUMB[16][5] ) );
  FAX1 S3_15_6 ( .A(n40), .B(\CARRYB[14][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[15][6] ), .YS(\SUMB[15][6] ) );
  FAX1 S2_15_5 ( .A(n39), .B(\CARRYB[14][5] ), .C(\SUMB[14][6] ), .YC(
        \CARRYB[15][5] ), .YS(\SUMB[15][5] ) );
  FAX1 S3_14_6 ( .A(n40), .B(\CARRYB[13][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[14][6] ), .YS(\SUMB[14][6] ) );
  FAX1 S2_14_5 ( .A(n39), .B(\CARRYB[13][5] ), .C(\SUMB[13][6] ), .YC(
        \CARRYB[14][5] ), .YS(\SUMB[14][5] ) );
  FAX1 S3_13_6 ( .A(n40), .B(\CARRYB[12][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[13][6] ), .YS(\SUMB[13][6] ) );
  FAX1 S2_13_5 ( .A(n39), .B(\CARRYB[12][5] ), .C(\SUMB[12][6] ), .YC(
        \CARRYB[13][5] ), .YS(\SUMB[13][5] ) );
  FAX1 S3_12_6 ( .A(n40), .B(\CARRYB[11][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[12][6] ), .YS(\SUMB[12][6] ) );
  FAX1 S2_12_5 ( .A(n39), .B(\CARRYB[11][5] ), .C(\SUMB[11][6] ), .YC(
        \CARRYB[12][5] ), .YS(\SUMB[12][5] ) );
  FAX1 S3_11_6 ( .A(n40), .B(\CARRYB[10][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[11][6] ), .YS(\SUMB[11][6] ) );
  FAX1 S2_11_5 ( .A(n39), .B(\CARRYB[10][5] ), .C(\SUMB[10][6] ), .YC(
        \CARRYB[11][5] ), .YS(\SUMB[11][5] ) );
  FAX1 S3_10_6 ( .A(n40), .B(\CARRYB[9][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[10][6] ), .YS(\SUMB[10][6] ) );
  FAX1 S2_10_5 ( .A(n39), .B(\CARRYB[9][5] ), .C(\SUMB[9][6] ), .YC(
        \CARRYB[10][5] ), .YS(\SUMB[10][5] ) );
  FAX1 S3_9_6 ( .A(n40), .B(\CARRYB[8][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[9][6] ), .YS(\SUMB[9][6] ) );
  FAX1 S2_9_5 ( .A(n39), .B(\CARRYB[8][5] ), .C(\SUMB[8][6] ), .YC(
        \CARRYB[9][5] ), .YS(\SUMB[9][5] ) );
  FAX1 S3_8_6 ( .A(n40), .B(\CARRYB[7][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[8][6] ), .YS(\SUMB[8][6] ) );
  FAX1 S2_8_5 ( .A(n39), .B(\CARRYB[7][5] ), .C(\SUMB[7][6] ), .YC(
        \CARRYB[8][5] ), .YS(\SUMB[8][5] ) );
  FAX1 S3_7_6 ( .A(n40), .B(\CARRYB[6][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S2_7_5 ( .A(n39), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S3_6_6 ( .A(n40), .B(\CARRYB[5][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_5 ( .A(n39), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S3_5_6 ( .A(n40), .B(\CARRYB[4][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_5 ( .A(n39), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S3_4_6 ( .A(n40), .B(\CARRYB[3][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_5 ( .A(n39), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S3_3_6 ( .A(n40), .B(\CARRYB[2][6] ), .C(\ab[9][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  AND2X2 U9 ( .A(B[7]), .B(A[9]), .Y(\ab[9][7] ) );
  FAX1 S2_3_5 ( .A(n39), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S3_2_6 ( .A(n40), .B(n4), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), .YS(
        \SUMB[2][6] ) );
  NAND2X1 U10 ( .A(B[6]), .B(A[9]), .Y(n10) );
  FAX1 S2_2_5 ( .A(n39), .B(n3), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), .YS(
        \SUMB[2][5] ) );
  NAND2X1 U12 ( .A(B[5]), .B(A[9]), .Y(n12) );
  INVX4 U11 ( .A(n10), .Y(n40) );
  INVX4 U13 ( .A(n12), .Y(n39) );
  INVX4 U15 ( .A(n14), .Y(n38) );
  INVX4 U17 ( .A(n16), .Y(n37) );
  INVX4 U19 ( .A(n18), .Y(n36) );
  INVX4 U21 ( .A(n20), .Y(n35) );
  INVX4 U23 ( .A(n22), .Y(n34) );
  INVX2 U31 ( .A(A[1]), .Y(n41) );
  INVX2 U32 ( .A(A[0]), .Y(n42) );
  INVX2 U33 ( .A(B[0]), .Y(n43) );
  INVX2 U34 ( .A(B[1]), .Y(n44) );
  INVX2 U35 ( .A(B[2]), .Y(n45) );
  INVX2 U36 ( .A(B[3]), .Y(n46) );
  INVX2 U37 ( .A(B[4]), .Y(n47) );
  INVX2 U38 ( .A(B[5]), .Y(n48) );
  INVX2 U39 ( .A(B[6]), .Y(n49) );
  INVX2 U40 ( .A(B[7]), .Y(n50) );
endmodule


module CannyEdge_DW02_mult_14 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] , n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n60, n61, n62;
  assign \ab[1][7]  = B[7];
  assign \ab[1][6]  = B[6];
  assign \ab[1][5]  = B[5];
  assign \ab[1][4]  = B[4];
  assign \ab[1][3]  = B[3];
  assign \ab[1][2]  = B[2];
  assign \ab[1][1]  = B[1];
  assign PRODUCT[0] = \ab[1][0] ;
  assign \ab[1][0]  = B[0];

  AND2X2 U2 ( .A(n35), .B(\SUMB[6][4] ), .Y(n3) );
  AND2X2 U3 ( .A(n32), .B(\SUMB[6][1] ), .Y(n4) );
  AND2X2 U4 ( .A(n36), .B(\SUMB[2][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n37), .B(\SUMB[2][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[2][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n39), .B(\SUMB[2][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n40), .B(\SUMB[2][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n41), .B(\SUMB[2][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n27), .B(\SUMB[4][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n33), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n34), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n11), .B(n43), .Y(n14) );
  AND2X2 U14 ( .A(\ab[1][2] ), .B(\ab[1][1] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[1][3] ), .B(\ab[1][2] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[1][4] ), .B(\ab[1][3] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[1][5] ), .B(\ab[1][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[1][6] ), .B(\ab[1][5] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[1][7] ), .B(\ab[1][6] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[1][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n4), .B(\SUMB[7][1] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[3][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[3][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[3][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[3][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][5] ), .Y(n27) );
  AND2X2 U27 ( .A(n23), .B(\SUMB[4][1] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[4][2] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[4][3] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[4][4] ), .Y(n31) );
  AND2X2 U31 ( .A(n28), .B(\SUMB[5][1] ), .Y(n32) );
  AND2X2 U32 ( .A(n29), .B(\SUMB[5][2] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][3] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][4] ), .Y(n35) );
  AND2X2 U35 ( .A(n21), .B(\SUMB[1][1] ), .Y(n36) );
  AND2X2 U36 ( .A(n15), .B(\SUMB[1][2] ), .Y(n37) );
  AND2X2 U37 ( .A(n16), .B(\SUMB[1][3] ), .Y(n38) );
  AND2X2 U38 ( .A(n17), .B(\SUMB[1][4] ), .Y(n39) );
  AND2X2 U39 ( .A(n18), .B(\SUMB[1][5] ), .Y(n40) );
  AND2X2 U40 ( .A(n19), .B(\SUMB[1][6] ), .Y(n41) );
  AND2X2 U41 ( .A(n20), .B(\ab[1][7] ), .Y(n42) );
  AND2X2 U42 ( .A(n10), .B(n42), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n13), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n12), .Y(n45) );
  XNOR2X1 U45 ( .A(n61), .B(n22), .Y(PRODUCT[9]) );
  XOR2X1 U46 ( .A(\SUMB[7][1] ), .B(n4), .Y(PRODUCT[8]) );
  XOR2X1 U47 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U48 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U49 ( .A(n14), .B(n3), .Y(\A1[9] ) );
  NAND2X1 U50 ( .A(n14), .B(n3), .Y(n47) );
  XOR2X1 U51 ( .A(\ab[1][0] ), .B(\ab[1][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U52 ( .A(\ab[1][1] ), .B(\ab[1][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U53 ( .A(\ab[1][2] ), .B(\ab[1][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U54 ( .A(\ab[1][3] ), .B(\ab[1][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U55 ( .A(\ab[1][4] ), .B(\ab[1][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U56 ( .A(\ab[1][5] ), .B(\ab[1][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U57 ( .A(\ab[1][6] ), .B(\ab[1][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U58 ( .A(\SUMB[1][1] ), .B(n21), .Y(PRODUCT[2]) );
  XOR2X1 U59 ( .A(\SUMB[1][2] ), .B(n15), .Y(\SUMB[2][1] ) );
  XOR2X1 U60 ( .A(\SUMB[1][3] ), .B(n16), .Y(\SUMB[2][2] ) );
  XOR2X1 U61 ( .A(\SUMB[1][4] ), .B(n17), .Y(\SUMB[2][3] ) );
  XOR2X1 U62 ( .A(\SUMB[1][5] ), .B(n18), .Y(\SUMB[2][4] ) );
  XOR2X1 U63 ( .A(\SUMB[1][6] ), .B(n19), .Y(\SUMB[2][5] ) );
  XOR2X1 U64 ( .A(\ab[1][7] ), .B(n20), .Y(\SUMB[2][6] ) );
  XOR2X1 U65 ( .A(\SUMB[2][1] ), .B(n36), .Y(PRODUCT[3]) );
  XOR2X1 U66 ( .A(\SUMB[2][2] ), .B(n37), .Y(\SUMB[3][1] ) );
  XOR2X1 U67 ( .A(\SUMB[2][3] ), .B(n38), .Y(\SUMB[3][2] ) );
  XOR2X1 U68 ( .A(\SUMB[2][4] ), .B(n39), .Y(\SUMB[3][3] ) );
  XOR2X1 U69 ( .A(\SUMB[2][5] ), .B(n40), .Y(\SUMB[3][4] ) );
  XOR2X1 U70 ( .A(\SUMB[2][6] ), .B(n41), .Y(\SUMB[3][5] ) );
  XOR2X1 U71 ( .A(\SUMB[3][1] ), .B(n5), .Y(PRODUCT[4]) );
  XOR2X1 U72 ( .A(\SUMB[3][2] ), .B(n6), .Y(\SUMB[4][1] ) );
  XOR2X1 U73 ( .A(\SUMB[3][3] ), .B(n7), .Y(\SUMB[4][2] ) );
  XOR2X1 U74 ( .A(\SUMB[3][4] ), .B(n8), .Y(\SUMB[4][3] ) );
  XOR2X1 U75 ( .A(\SUMB[3][5] ), .B(n9), .Y(\SUMB[4][4] ) );
  XOR2X1 U76 ( .A(n42), .B(n10), .Y(\SUMB[4][5] ) );
  XOR2X1 U77 ( .A(\SUMB[4][1] ), .B(n23), .Y(PRODUCT[5]) );
  XOR2X1 U78 ( .A(\SUMB[4][2] ), .B(n24), .Y(\SUMB[5][1] ) );
  XOR2X1 U79 ( .A(\SUMB[4][3] ), .B(n25), .Y(\SUMB[5][2] ) );
  XOR2X1 U80 ( .A(\SUMB[4][4] ), .B(n26), .Y(\SUMB[5][3] ) );
  XOR2X1 U81 ( .A(\SUMB[4][5] ), .B(n27), .Y(\SUMB[5][4] ) );
  XOR2X1 U82 ( .A(\SUMB[5][1] ), .B(n28), .Y(PRODUCT[6]) );
  XOR2X1 U83 ( .A(\SUMB[5][2] ), .B(n29), .Y(\SUMB[6][1] ) );
  XOR2X1 U84 ( .A(\SUMB[5][3] ), .B(n30), .Y(\SUMB[6][2] ) );
  XOR2X1 U85 ( .A(\SUMB[5][4] ), .B(n31), .Y(\SUMB[6][3] ) );
  XOR2X1 U86 ( .A(n43), .B(n11), .Y(\SUMB[6][4] ) );
  XOR2X1 U87 ( .A(\SUMB[6][1] ), .B(n32), .Y(PRODUCT[7]) );
  XOR2X1 U88 ( .A(\SUMB[6][2] ), .B(n33), .Y(\SUMB[7][1] ) );
  XOR2X1 U89 ( .A(\SUMB[6][3] ), .B(n34), .Y(\SUMB[7][2] ) );
  XOR2X1 U90 ( .A(\SUMB[6][4] ), .B(n35), .Y(\SUMB[7][3] ) );
  NOR2X1 U91 ( .A(n45), .B(\A1[8] ), .Y(n50) );
  NAND2X1 U92 ( .A(n45), .B(\A1[8] ), .Y(n51) );
  OAI21X1 U93 ( .A(n48), .B(n50), .C(n51), .Y(n56) );
  NOR2X1 U94 ( .A(n44), .B(\A1[9] ), .Y(n53) );
  AND2X1 U95 ( .A(n44), .B(\A1[9] ), .Y(n54) );
  AOI21X1 U96 ( .A(n56), .B(n62), .C(n54), .Y(n49) );
  XOR2X1 U97 ( .A(n47), .B(n49), .Y(PRODUCT[12]) );
  NAND2X1 U98 ( .A(n60), .B(n51), .Y(n52) );
  XOR2X1 U99 ( .A(n52), .B(n48), .Y(PRODUCT[10]) );
  NOR2X1 U100 ( .A(n54), .B(n53), .Y(n55) );
  XOR2X1 U101 ( .A(n56), .B(n55), .Y(PRODUCT[11]) );
  NAND2X1 U102 ( .A(\A1[7] ), .B(n22), .Y(n48) );
  NOR2X1 U103 ( .A(n47), .B(n49), .Y(PRODUCT[13]) );
  INVX2 U104 ( .A(n50), .Y(n60) );
  INVX2 U105 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U106 ( .A(n53), .Y(n62) );
endmodule


module CannyEdge_DW02_mult_15 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [7:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , n9, n8, n7, n6, n5, n4, n3, n24, n22, n20,
         n18, n16, n14, n12, n10, \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[30][1] ,
         \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] ,
         \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[30][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] ,
         \CARRYB[28][1] , \CARRYB[28][0] , \CARRYB[27][3] , \CARRYB[27][2] ,
         \CARRYB[27][1] , \CARRYB[27][0] , \CARRYB[26][4] , \CARRYB[26][3] ,
         \CARRYB[26][2] , \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] ,
         \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][6] ,
         \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] ,
         \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][6] ,
         \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] ,
         \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] ,
         \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][6] ,
         \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] ,
         \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , n26, n27, n28, n29, n30, n31, n32,
         n33;

  XOR2X1 U31 ( .A(n33), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  AND2X1 U32 ( .A(B[7]), .B(A[0]), .Y(\ab[0][7] ) );
  AND2X1 U33 ( .A(B[6]), .B(A[0]), .Y(\ab[0][6] ) );
  AND2X1 U34 ( .A(B[5]), .B(A[0]), .Y(\ab[0][5] ) );
  AND2X1 U35 ( .A(B[4]), .B(A[0]), .Y(\ab[0][4] ) );
  AND2X1 U36 ( .A(B[3]), .B(A[0]), .Y(\ab[0][3] ) );
  AND2X1 U37 ( .A(B[2]), .B(A[0]), .Y(\ab[0][2] ) );
  AND2X1 U38 ( .A(B[1]), .B(A[0]), .Y(\ab[0][1] ) );
  AND2X1 U39 ( .A(B[0]), .B(A[0]), .Y(PRODUCT[0]) );
  FAX1 S4_0 ( .A(n33), .B(\CARRYB[30][0] ), .C(\SUMB[30][1] ), .YS(PRODUCT[31]) );
  FAX1 S1_30_0 ( .A(n33), .B(\CARRYB[29][0] ), .C(\SUMB[29][1] ), .YC(
        \CARRYB[30][0] ), .YS(PRODUCT[30]) );
  FAX1 S1_29_0 ( .A(n33), .B(\CARRYB[28][0] ), .C(\SUMB[28][1] ), .YC(
        \CARRYB[29][0] ), .YS(PRODUCT[29]) );
  FAX1 S1_28_0 ( .A(n33), .B(\CARRYB[27][0] ), .C(\SUMB[27][1] ), .YC(
        \CARRYB[28][0] ), .YS(PRODUCT[28]) );
  FAX1 S1_27_0 ( .A(n33), .B(\CARRYB[26][0] ), .C(\SUMB[26][1] ), .YC(
        \CARRYB[27][0] ), .YS(PRODUCT[27]) );
  FAX1 S1_26_0 ( .A(n33), .B(\CARRYB[25][0] ), .C(\SUMB[25][1] ), .YC(
        \CARRYB[26][0] ), .YS(PRODUCT[26]) );
  FAX1 S1_25_0 ( .A(n33), .B(\CARRYB[24][0] ), .C(\SUMB[24][1] ), .YC(
        \CARRYB[25][0] ), .YS(PRODUCT[25]) );
  FAX1 S1_24_0 ( .A(n33), .B(\CARRYB[23][0] ), .C(\SUMB[23][1] ), .YC(
        \CARRYB[24][0] ), .YS(PRODUCT[24]) );
  FAX1 S1_23_0 ( .A(n33), .B(\CARRYB[22][0] ), .C(\SUMB[22][1] ), .YC(
        \CARRYB[23][0] ), .YS(PRODUCT[23]) );
  FAX1 S1_22_0 ( .A(n33), .B(\CARRYB[21][0] ), .C(\SUMB[21][1] ), .YC(
        \CARRYB[22][0] ), .YS(PRODUCT[22]) );
  FAX1 S1_21_0 ( .A(n33), .B(\CARRYB[20][0] ), .C(\SUMB[20][1] ), .YC(
        \CARRYB[21][0] ), .YS(PRODUCT[21]) );
  FAX1 S1_20_0 ( .A(n33), .B(\CARRYB[19][0] ), .C(\SUMB[19][1] ), .YC(
        \CARRYB[20][0] ), .YS(PRODUCT[20]) );
  FAX1 S1_19_0 ( .A(n33), .B(\CARRYB[18][0] ), .C(\SUMB[18][1] ), .YC(
        \CARRYB[19][0] ), .YS(PRODUCT[19]) );
  FAX1 S1_18_0 ( .A(n33), .B(\CARRYB[17][0] ), .C(\SUMB[17][1] ), .YC(
        \CARRYB[18][0] ), .YS(PRODUCT[18]) );
  FAX1 S1_17_0 ( .A(n33), .B(\CARRYB[16][0] ), .C(\SUMB[16][1] ), .YC(
        \CARRYB[17][0] ), .YS(PRODUCT[17]) );
  FAX1 S1_16_0 ( .A(n33), .B(\CARRYB[15][0] ), .C(\SUMB[15][1] ), .YC(
        \CARRYB[16][0] ), .YS(PRODUCT[16]) );
  FAX1 S1_15_0 ( .A(n33), .B(\CARRYB[14][0] ), .C(\SUMB[14][1] ), .YC(
        \CARRYB[15][0] ), .YS(PRODUCT[15]) );
  FAX1 S1_14_0 ( .A(n33), .B(\CARRYB[13][0] ), .C(\SUMB[13][1] ), .YC(
        \CARRYB[14][0] ), .YS(PRODUCT[14]) );
  FAX1 S1_13_0 ( .A(n33), .B(\CARRYB[12][0] ), .C(\SUMB[12][1] ), .YC(
        \CARRYB[13][0] ), .YS(PRODUCT[13]) );
  FAX1 S1_12_0 ( .A(n33), .B(\CARRYB[11][0] ), .C(\SUMB[11][1] ), .YC(
        \CARRYB[12][0] ), .YS(PRODUCT[12]) );
  FAX1 S1_11_0 ( .A(n33), .B(\CARRYB[10][0] ), .C(\SUMB[10][1] ), .YC(
        \CARRYB[11][0] ), .YS(PRODUCT[11]) );
  FAX1 S1_10_0 ( .A(n33), .B(\CARRYB[9][0] ), .C(\SUMB[9][1] ), .YC(
        \CARRYB[10][0] ), .YS(PRODUCT[10]) );
  FAX1 S1_9_0 ( .A(n33), .B(\CARRYB[8][0] ), .C(\SUMB[8][1] ), .YC(
        \CARRYB[9][0] ), .YS(PRODUCT[9]) );
  FAX1 S1_8_0 ( .A(n33), .B(\CARRYB[7][0] ), .C(\SUMB[7][1] ), .YC(
        \CARRYB[8][0] ), .YS(PRODUCT[8]) );
  FAX1 S1_7_0 ( .A(n33), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(PRODUCT[7]) );
  FAX1 S1_6_0 ( .A(n33), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(PRODUCT[6]) );
  FAX1 S1_5_0 ( .A(n33), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(PRODUCT[5]) );
  FAX1 S1_4_0 ( .A(n33), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(PRODUCT[4]) );
  FAX1 S1_3_0 ( .A(n33), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(PRODUCT[3]) );
  FAX1 S1_2_0 ( .A(n33), .B(n3), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), .YS(
        PRODUCT[2]) );
  XOR2X1 U30 ( .A(n26), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  AND2X2 U2 ( .A(\ab[0][1] ), .B(n33), .Y(n3) );
  NAND2X1 U23 ( .A(B[0]), .B(A[9]), .Y(n24) );
  FAX1 S2_30_1 ( .A(n26), .B(\CARRYB[29][1] ), .C(\SUMB[29][2] ), .YS(
        \SUMB[30][1] ) );
  FAX1 S2_29_1 ( .A(n26), .B(\CARRYB[28][1] ), .C(\SUMB[28][2] ), .YC(
        \CARRYB[29][1] ), .YS(\SUMB[29][1] ) );
  FAX1 S2_28_1 ( .A(n26), .B(\CARRYB[27][1] ), .C(\SUMB[27][2] ), .YC(
        \CARRYB[28][1] ), .YS(\SUMB[28][1] ) );
  FAX1 S2_27_1 ( .A(n26), .B(\CARRYB[26][1] ), .C(\SUMB[26][2] ), .YC(
        \CARRYB[27][1] ), .YS(\SUMB[27][1] ) );
  FAX1 S2_26_1 ( .A(n26), .B(\CARRYB[25][1] ), .C(\SUMB[25][2] ), .YC(
        \CARRYB[26][1] ), .YS(\SUMB[26][1] ) );
  FAX1 S2_25_1 ( .A(n26), .B(\CARRYB[24][1] ), .C(\SUMB[24][2] ), .YC(
        \CARRYB[25][1] ), .YS(\SUMB[25][1] ) );
  FAX1 S2_24_1 ( .A(n26), .B(\CARRYB[23][1] ), .C(\SUMB[23][2] ), .YC(
        \CARRYB[24][1] ), .YS(\SUMB[24][1] ) );
  FAX1 S2_23_1 ( .A(n26), .B(\CARRYB[22][1] ), .C(\SUMB[22][2] ), .YC(
        \CARRYB[23][1] ), .YS(\SUMB[23][1] ) );
  FAX1 S2_22_1 ( .A(n26), .B(\CARRYB[21][1] ), .C(\SUMB[21][2] ), .YC(
        \CARRYB[22][1] ), .YS(\SUMB[22][1] ) );
  FAX1 S2_21_1 ( .A(n26), .B(\CARRYB[20][1] ), .C(\SUMB[20][2] ), .YC(
        \CARRYB[21][1] ), .YS(\SUMB[21][1] ) );
  FAX1 S2_20_1 ( .A(n26), .B(\CARRYB[19][1] ), .C(\SUMB[19][2] ), .YC(
        \CARRYB[20][1] ), .YS(\SUMB[20][1] ) );
  FAX1 S2_19_1 ( .A(n26), .B(\CARRYB[18][1] ), .C(\SUMB[18][2] ), .YC(
        \CARRYB[19][1] ), .YS(\SUMB[19][1] ) );
  FAX1 S2_18_1 ( .A(n26), .B(\CARRYB[17][1] ), .C(\SUMB[17][2] ), .YC(
        \CARRYB[18][1] ), .YS(\SUMB[18][1] ) );
  FAX1 S2_17_1 ( .A(n26), .B(\CARRYB[16][1] ), .C(\SUMB[16][2] ), .YC(
        \CARRYB[17][1] ), .YS(\SUMB[17][1] ) );
  FAX1 S2_16_1 ( .A(n26), .B(\CARRYB[15][1] ), .C(\SUMB[15][2] ), .YC(
        \CARRYB[16][1] ), .YS(\SUMB[16][1] ) );
  FAX1 S2_15_1 ( .A(n26), .B(\CARRYB[14][1] ), .C(\SUMB[14][2] ), .YC(
        \CARRYB[15][1] ), .YS(\SUMB[15][1] ) );
  FAX1 S2_14_1 ( .A(n26), .B(\CARRYB[13][1] ), .C(\SUMB[13][2] ), .YC(
        \CARRYB[14][1] ), .YS(\SUMB[14][1] ) );
  FAX1 S2_13_1 ( .A(n26), .B(\CARRYB[12][1] ), .C(\SUMB[12][2] ), .YC(
        \CARRYB[13][1] ), .YS(\SUMB[13][1] ) );
  FAX1 S2_12_1 ( .A(n26), .B(\CARRYB[11][1] ), .C(\SUMB[11][2] ), .YC(
        \CARRYB[12][1] ), .YS(\SUMB[12][1] ) );
  FAX1 S2_11_1 ( .A(n26), .B(\CARRYB[10][1] ), .C(\SUMB[10][2] ), .YC(
        \CARRYB[11][1] ), .YS(\SUMB[11][1] ) );
  FAX1 S2_10_1 ( .A(n26), .B(\CARRYB[9][1] ), .C(\SUMB[9][2] ), .YC(
        \CARRYB[10][1] ), .YS(\SUMB[10][1] ) );
  FAX1 S2_9_1 ( .A(n26), .B(\CARRYB[8][1] ), .C(\SUMB[8][2] ), .YC(
        \CARRYB[9][1] ), .YS(\SUMB[9][1] ) );
  FAX1 S2_8_1 ( .A(n26), .B(\CARRYB[7][1] ), .C(\SUMB[7][2] ), .YC(
        \CARRYB[8][1] ), .YS(\SUMB[8][1] ) );
  FAX1 S2_7_1 ( .A(n26), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S2_6_1 ( .A(n26), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_5_1 ( .A(n26), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_4_1 ( .A(n26), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_3_1 ( .A(n26), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_2_1 ( .A(n26), .B(n4), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), .YS(
        \SUMB[2][1] ) );
  XOR2X1 U29 ( .A(n27), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  AND2X2 U3 ( .A(\ab[0][2] ), .B(n26), .Y(n4) );
  NAND2X1 U21 ( .A(B[1]), .B(A[9]), .Y(n22) );
  FAX1 S2_29_2 ( .A(n27), .B(\CARRYB[28][2] ), .C(\SUMB[28][3] ), .YS(
        \SUMB[29][2] ) );
  FAX1 S2_28_2 ( .A(n27), .B(\CARRYB[27][2] ), .C(\SUMB[27][3] ), .YC(
        \CARRYB[28][2] ), .YS(\SUMB[28][2] ) );
  FAX1 S2_27_2 ( .A(n27), .B(\CARRYB[26][2] ), .C(\SUMB[26][3] ), .YC(
        \CARRYB[27][2] ), .YS(\SUMB[27][2] ) );
  FAX1 S2_26_2 ( .A(n27), .B(\CARRYB[25][2] ), .C(\SUMB[25][3] ), .YC(
        \CARRYB[26][2] ), .YS(\SUMB[26][2] ) );
  FAX1 S2_25_2 ( .A(n27), .B(\CARRYB[24][2] ), .C(\SUMB[24][3] ), .YC(
        \CARRYB[25][2] ), .YS(\SUMB[25][2] ) );
  FAX1 S2_24_2 ( .A(n27), .B(\CARRYB[23][2] ), .C(\SUMB[23][3] ), .YC(
        \CARRYB[24][2] ), .YS(\SUMB[24][2] ) );
  FAX1 S2_23_2 ( .A(n27), .B(\CARRYB[22][2] ), .C(\SUMB[22][3] ), .YC(
        \CARRYB[23][2] ), .YS(\SUMB[23][2] ) );
  FAX1 S2_22_2 ( .A(n27), .B(\CARRYB[21][2] ), .C(\SUMB[21][3] ), .YC(
        \CARRYB[22][2] ), .YS(\SUMB[22][2] ) );
  FAX1 S2_21_2 ( .A(n27), .B(\CARRYB[20][2] ), .C(\SUMB[20][3] ), .YC(
        \CARRYB[21][2] ), .YS(\SUMB[21][2] ) );
  FAX1 S2_20_2 ( .A(n27), .B(\CARRYB[19][2] ), .C(\SUMB[19][3] ), .YC(
        \CARRYB[20][2] ), .YS(\SUMB[20][2] ) );
  FAX1 S2_19_2 ( .A(n27), .B(\CARRYB[18][2] ), .C(\SUMB[18][3] ), .YC(
        \CARRYB[19][2] ), .YS(\SUMB[19][2] ) );
  FAX1 S2_18_2 ( .A(n27), .B(\CARRYB[17][2] ), .C(\SUMB[17][3] ), .YC(
        \CARRYB[18][2] ), .YS(\SUMB[18][2] ) );
  FAX1 S2_17_2 ( .A(n27), .B(\CARRYB[16][2] ), .C(\SUMB[16][3] ), .YC(
        \CARRYB[17][2] ), .YS(\SUMB[17][2] ) );
  FAX1 S2_16_2 ( .A(n27), .B(\CARRYB[15][2] ), .C(\SUMB[15][3] ), .YC(
        \CARRYB[16][2] ), .YS(\SUMB[16][2] ) );
  FAX1 S2_15_2 ( .A(n27), .B(\CARRYB[14][2] ), .C(\SUMB[14][3] ), .YC(
        \CARRYB[15][2] ), .YS(\SUMB[15][2] ) );
  FAX1 S2_14_2 ( .A(n27), .B(\CARRYB[13][2] ), .C(\SUMB[13][3] ), .YC(
        \CARRYB[14][2] ), .YS(\SUMB[14][2] ) );
  FAX1 S2_13_2 ( .A(n27), .B(\CARRYB[12][2] ), .C(\SUMB[12][3] ), .YC(
        \CARRYB[13][2] ), .YS(\SUMB[13][2] ) );
  FAX1 S2_12_2 ( .A(n27), .B(\CARRYB[11][2] ), .C(\SUMB[11][3] ), .YC(
        \CARRYB[12][2] ), .YS(\SUMB[12][2] ) );
  FAX1 S2_11_2 ( .A(n27), .B(\CARRYB[10][2] ), .C(\SUMB[10][3] ), .YC(
        \CARRYB[11][2] ), .YS(\SUMB[11][2] ) );
  FAX1 S2_10_2 ( .A(n27), .B(\CARRYB[9][2] ), .C(\SUMB[9][3] ), .YC(
        \CARRYB[10][2] ), .YS(\SUMB[10][2] ) );
  FAX1 S2_9_2 ( .A(n27), .B(\CARRYB[8][2] ), .C(\SUMB[8][3] ), .YC(
        \CARRYB[9][2] ), .YS(\SUMB[9][2] ) );
  FAX1 S2_8_2 ( .A(n27), .B(\CARRYB[7][2] ), .C(\SUMB[7][3] ), .YC(
        \CARRYB[8][2] ), .YS(\SUMB[8][2] ) );
  FAX1 S2_7_2 ( .A(n27), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(n27), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_5_2 ( .A(n27), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_4_2 ( .A(n27), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_3_2 ( .A(n27), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_2_2 ( .A(n27), .B(n5), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), .YS(
        \SUMB[2][2] ) );
  XOR2X1 U28 ( .A(n29), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  AND2X2 U4 ( .A(\ab[0][3] ), .B(n27), .Y(n5) );
  NAND2X1 U19 ( .A(B[2]), .B(A[9]), .Y(n20) );
  FAX1 S2_28_3 ( .A(n29), .B(\CARRYB[27][3] ), .C(\SUMB[27][4] ), .YS(
        \SUMB[28][3] ) );
  FAX1 S2_27_3 ( .A(n29), .B(\CARRYB[26][3] ), .C(\SUMB[26][4] ), .YC(
        \CARRYB[27][3] ), .YS(\SUMB[27][3] ) );
  FAX1 S2_26_3 ( .A(n29), .B(\CARRYB[25][3] ), .C(\SUMB[25][4] ), .YC(
        \CARRYB[26][3] ), .YS(\SUMB[26][3] ) );
  FAX1 S2_25_3 ( .A(n29), .B(\CARRYB[24][3] ), .C(\SUMB[24][4] ), .YC(
        \CARRYB[25][3] ), .YS(\SUMB[25][3] ) );
  FAX1 S2_24_3 ( .A(n29), .B(\CARRYB[23][3] ), .C(\SUMB[23][4] ), .YC(
        \CARRYB[24][3] ), .YS(\SUMB[24][3] ) );
  FAX1 S2_23_3 ( .A(n29), .B(\CARRYB[22][3] ), .C(\SUMB[22][4] ), .YC(
        \CARRYB[23][3] ), .YS(\SUMB[23][3] ) );
  FAX1 S2_22_3 ( .A(n29), .B(\CARRYB[21][3] ), .C(\SUMB[21][4] ), .YC(
        \CARRYB[22][3] ), .YS(\SUMB[22][3] ) );
  FAX1 S2_21_3 ( .A(n29), .B(\CARRYB[20][3] ), .C(\SUMB[20][4] ), .YC(
        \CARRYB[21][3] ), .YS(\SUMB[21][3] ) );
  FAX1 S2_20_3 ( .A(n29), .B(\CARRYB[19][3] ), .C(\SUMB[19][4] ), .YC(
        \CARRYB[20][3] ), .YS(\SUMB[20][3] ) );
  FAX1 S2_19_3 ( .A(n29), .B(\CARRYB[18][3] ), .C(\SUMB[18][4] ), .YC(
        \CARRYB[19][3] ), .YS(\SUMB[19][3] ) );
  FAX1 S2_18_3 ( .A(n29), .B(\CARRYB[17][3] ), .C(\SUMB[17][4] ), .YC(
        \CARRYB[18][3] ), .YS(\SUMB[18][3] ) );
  FAX1 S2_17_3 ( .A(n29), .B(\CARRYB[16][3] ), .C(\SUMB[16][4] ), .YC(
        \CARRYB[17][3] ), .YS(\SUMB[17][3] ) );
  FAX1 S2_16_3 ( .A(n29), .B(\CARRYB[15][3] ), .C(\SUMB[15][4] ), .YC(
        \CARRYB[16][3] ), .YS(\SUMB[16][3] ) );
  FAX1 S2_15_3 ( .A(n29), .B(\CARRYB[14][3] ), .C(\SUMB[14][4] ), .YC(
        \CARRYB[15][3] ), .YS(\SUMB[15][3] ) );
  FAX1 S2_14_3 ( .A(n29), .B(\CARRYB[13][3] ), .C(\SUMB[13][4] ), .YC(
        \CARRYB[14][3] ), .YS(\SUMB[14][3] ) );
  FAX1 S2_13_3 ( .A(n29), .B(\CARRYB[12][3] ), .C(\SUMB[12][4] ), .YC(
        \CARRYB[13][3] ), .YS(\SUMB[13][3] ) );
  FAX1 S2_12_3 ( .A(n29), .B(\CARRYB[11][3] ), .C(\SUMB[11][4] ), .YC(
        \CARRYB[12][3] ), .YS(\SUMB[12][3] ) );
  FAX1 S2_11_3 ( .A(n29), .B(\CARRYB[10][3] ), .C(\SUMB[10][4] ), .YC(
        \CARRYB[11][3] ), .YS(\SUMB[11][3] ) );
  FAX1 S2_10_3 ( .A(n29), .B(\CARRYB[9][3] ), .C(\SUMB[9][4] ), .YC(
        \CARRYB[10][3] ), .YS(\SUMB[10][3] ) );
  FAX1 S2_9_3 ( .A(n29), .B(\CARRYB[8][3] ), .C(\SUMB[8][4] ), .YC(
        \CARRYB[9][3] ), .YS(\SUMB[9][3] ) );
  FAX1 S2_8_3 ( .A(n29), .B(\CARRYB[7][3] ), .C(\SUMB[7][4] ), .YC(
        \CARRYB[8][3] ), .YS(\SUMB[8][3] ) );
  FAX1 S2_7_3 ( .A(n29), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(n29), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(n29), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_4_3 ( .A(n29), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_3_3 ( .A(n29), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_2_3 ( .A(n29), .B(n6), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), .YS(
        \SUMB[2][3] ) );
  XOR2X1 U27 ( .A(n28), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  AND2X2 U5 ( .A(\ab[0][4] ), .B(n29), .Y(n6) );
  NAND2X1 U15 ( .A(B[3]), .B(A[9]), .Y(n16) );
  FAX1 S2_27_4 ( .A(n28), .B(\CARRYB[26][4] ), .C(\SUMB[26][5] ), .YS(
        \SUMB[27][4] ) );
  FAX1 S2_26_4 ( .A(n28), .B(\CARRYB[25][4] ), .C(\SUMB[25][5] ), .YC(
        \CARRYB[26][4] ), .YS(\SUMB[26][4] ) );
  FAX1 S2_25_4 ( .A(n28), .B(\CARRYB[24][4] ), .C(\SUMB[24][5] ), .YC(
        \CARRYB[25][4] ), .YS(\SUMB[25][4] ) );
  FAX1 S2_24_4 ( .A(n28), .B(\CARRYB[23][4] ), .C(\SUMB[23][5] ), .YC(
        \CARRYB[24][4] ), .YS(\SUMB[24][4] ) );
  FAX1 S2_23_4 ( .A(n28), .B(\CARRYB[22][4] ), .C(\SUMB[22][5] ), .YC(
        \CARRYB[23][4] ), .YS(\SUMB[23][4] ) );
  FAX1 S2_22_4 ( .A(n28), .B(\CARRYB[21][4] ), .C(\SUMB[21][5] ), .YC(
        \CARRYB[22][4] ), .YS(\SUMB[22][4] ) );
  FAX1 S2_21_4 ( .A(n28), .B(\CARRYB[20][4] ), .C(\SUMB[20][5] ), .YC(
        \CARRYB[21][4] ), .YS(\SUMB[21][4] ) );
  FAX1 S2_20_4 ( .A(n28), .B(\CARRYB[19][4] ), .C(\SUMB[19][5] ), .YC(
        \CARRYB[20][4] ), .YS(\SUMB[20][4] ) );
  FAX1 S2_19_4 ( .A(n28), .B(\CARRYB[18][4] ), .C(\SUMB[18][5] ), .YC(
        \CARRYB[19][4] ), .YS(\SUMB[19][4] ) );
  FAX1 S2_18_4 ( .A(n28), .B(\CARRYB[17][4] ), .C(\SUMB[17][5] ), .YC(
        \CARRYB[18][4] ), .YS(\SUMB[18][4] ) );
  FAX1 S2_17_4 ( .A(n28), .B(\CARRYB[16][4] ), .C(\SUMB[16][5] ), .YC(
        \CARRYB[17][4] ), .YS(\SUMB[17][4] ) );
  FAX1 S2_16_4 ( .A(n28), .B(\CARRYB[15][4] ), .C(\SUMB[15][5] ), .YC(
        \CARRYB[16][4] ), .YS(\SUMB[16][4] ) );
  FAX1 S2_15_4 ( .A(n28), .B(\CARRYB[14][4] ), .C(\SUMB[14][5] ), .YC(
        \CARRYB[15][4] ), .YS(\SUMB[15][4] ) );
  FAX1 S2_14_4 ( .A(n28), .B(\CARRYB[13][4] ), .C(\SUMB[13][5] ), .YC(
        \CARRYB[14][4] ), .YS(\SUMB[14][4] ) );
  FAX1 S2_13_4 ( .A(n28), .B(\CARRYB[12][4] ), .C(\SUMB[12][5] ), .YC(
        \CARRYB[13][4] ), .YS(\SUMB[13][4] ) );
  FAX1 S2_12_4 ( .A(n28), .B(\CARRYB[11][4] ), .C(\SUMB[11][5] ), .YC(
        \CARRYB[12][4] ), .YS(\SUMB[12][4] ) );
  FAX1 S2_11_4 ( .A(n28), .B(\CARRYB[10][4] ), .C(\SUMB[10][5] ), .YC(
        \CARRYB[11][4] ), .YS(\SUMB[11][4] ) );
  FAX1 S2_10_4 ( .A(n28), .B(\CARRYB[9][4] ), .C(\SUMB[9][5] ), .YC(
        \CARRYB[10][4] ), .YS(\SUMB[10][4] ) );
  FAX1 S2_9_4 ( .A(n28), .B(\CARRYB[8][4] ), .C(\SUMB[8][5] ), .YC(
        \CARRYB[9][4] ), .YS(\SUMB[9][4] ) );
  FAX1 S2_8_4 ( .A(n28), .B(\CARRYB[7][4] ), .C(\SUMB[7][5] ), .YC(
        \CARRYB[8][4] ), .YS(\SUMB[8][4] ) );
  FAX1 S2_7_4 ( .A(n28), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(n28), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(n28), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(n28), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_3_4 ( .A(n28), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_2_4 ( .A(n28), .B(n7), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), .YS(
        \SUMB[2][4] ) );
  XOR2X1 U26 ( .A(n30), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  AND2X2 U6 ( .A(\ab[0][5] ), .B(n28), .Y(n7) );
  NAND2X1 U17 ( .A(B[4]), .B(A[9]), .Y(n18) );
  FAX1 S2_26_5 ( .A(n30), .B(\CARRYB[25][5] ), .C(\SUMB[25][6] ), .YS(
        \SUMB[26][5] ) );
  FAX1 S3_25_6 ( .A(n31), .B(\CARRYB[24][6] ), .C(n32), .YS(\SUMB[25][6] ) );
  FAX1 S2_25_5 ( .A(n30), .B(\CARRYB[24][5] ), .C(\SUMB[24][6] ), .YC(
        \CARRYB[25][5] ), .YS(\SUMB[25][5] ) );
  FAX1 S3_24_6 ( .A(n31), .B(\CARRYB[23][6] ), .C(n32), .YC(\CARRYB[24][6] ), 
        .YS(\SUMB[24][6] ) );
  FAX1 S2_24_5 ( .A(n30), .B(\CARRYB[23][5] ), .C(\SUMB[23][6] ), .YC(
        \CARRYB[24][5] ), .YS(\SUMB[24][5] ) );
  FAX1 S3_23_6 ( .A(n31), .B(\CARRYB[22][6] ), .C(n32), .YC(\CARRYB[23][6] ), 
        .YS(\SUMB[23][6] ) );
  FAX1 S2_23_5 ( .A(n30), .B(\CARRYB[22][5] ), .C(\SUMB[22][6] ), .YC(
        \CARRYB[23][5] ), .YS(\SUMB[23][5] ) );
  FAX1 S3_22_6 ( .A(n31), .B(\CARRYB[21][6] ), .C(n32), .YC(\CARRYB[22][6] ), 
        .YS(\SUMB[22][6] ) );
  FAX1 S2_22_5 ( .A(n30), .B(\CARRYB[21][5] ), .C(\SUMB[21][6] ), .YC(
        \CARRYB[22][5] ), .YS(\SUMB[22][5] ) );
  FAX1 S3_21_6 ( .A(n31), .B(\CARRYB[20][6] ), .C(n32), .YC(\CARRYB[21][6] ), 
        .YS(\SUMB[21][6] ) );
  FAX1 S2_21_5 ( .A(n30), .B(\CARRYB[20][5] ), .C(\SUMB[20][6] ), .YC(
        \CARRYB[21][5] ), .YS(\SUMB[21][5] ) );
  FAX1 S3_20_6 ( .A(n31), .B(\CARRYB[19][6] ), .C(n32), .YC(\CARRYB[20][6] ), 
        .YS(\SUMB[20][6] ) );
  FAX1 S2_20_5 ( .A(n30), .B(\CARRYB[19][5] ), .C(\SUMB[19][6] ), .YC(
        \CARRYB[20][5] ), .YS(\SUMB[20][5] ) );
  FAX1 S3_19_6 ( .A(n31), .B(\CARRYB[18][6] ), .C(n32), .YC(\CARRYB[19][6] ), 
        .YS(\SUMB[19][6] ) );
  FAX1 S2_19_5 ( .A(n30), .B(\CARRYB[18][5] ), .C(\SUMB[18][6] ), .YC(
        \CARRYB[19][5] ), .YS(\SUMB[19][5] ) );
  FAX1 S3_18_6 ( .A(n31), .B(\CARRYB[17][6] ), .C(n32), .YC(\CARRYB[18][6] ), 
        .YS(\SUMB[18][6] ) );
  FAX1 S2_18_5 ( .A(n30), .B(\CARRYB[17][5] ), .C(\SUMB[17][6] ), .YC(
        \CARRYB[18][5] ), .YS(\SUMB[18][5] ) );
  FAX1 S3_17_6 ( .A(n31), .B(\CARRYB[16][6] ), .C(n32), .YC(\CARRYB[17][6] ), 
        .YS(\SUMB[17][6] ) );
  FAX1 S2_17_5 ( .A(n30), .B(\CARRYB[16][5] ), .C(\SUMB[16][6] ), .YC(
        \CARRYB[17][5] ), .YS(\SUMB[17][5] ) );
  FAX1 S3_16_6 ( .A(n31), .B(\CARRYB[15][6] ), .C(n32), .YC(\CARRYB[16][6] ), 
        .YS(\SUMB[16][6] ) );
  FAX1 S2_16_5 ( .A(n30), .B(\CARRYB[15][5] ), .C(\SUMB[15][6] ), .YC(
        \CARRYB[16][5] ), .YS(\SUMB[16][5] ) );
  FAX1 S3_15_6 ( .A(n31), .B(\CARRYB[14][6] ), .C(n32), .YC(\CARRYB[15][6] ), 
        .YS(\SUMB[15][6] ) );
  FAX1 S2_15_5 ( .A(n30), .B(\CARRYB[14][5] ), .C(\SUMB[14][6] ), .YC(
        \CARRYB[15][5] ), .YS(\SUMB[15][5] ) );
  FAX1 S3_14_6 ( .A(n31), .B(\CARRYB[13][6] ), .C(n32), .YC(\CARRYB[14][6] ), 
        .YS(\SUMB[14][6] ) );
  FAX1 S2_14_5 ( .A(n30), .B(\CARRYB[13][5] ), .C(\SUMB[13][6] ), .YC(
        \CARRYB[14][5] ), .YS(\SUMB[14][5] ) );
  FAX1 S3_13_6 ( .A(n31), .B(\CARRYB[12][6] ), .C(n32), .YC(\CARRYB[13][6] ), 
        .YS(\SUMB[13][6] ) );
  FAX1 S2_13_5 ( .A(n30), .B(\CARRYB[12][5] ), .C(\SUMB[12][6] ), .YC(
        \CARRYB[13][5] ), .YS(\SUMB[13][5] ) );
  FAX1 S3_12_6 ( .A(n31), .B(\CARRYB[11][6] ), .C(n32), .YC(\CARRYB[12][6] ), 
        .YS(\SUMB[12][6] ) );
  FAX1 S2_12_5 ( .A(n30), .B(\CARRYB[11][5] ), .C(\SUMB[11][6] ), .YC(
        \CARRYB[12][5] ), .YS(\SUMB[12][5] ) );
  FAX1 S3_11_6 ( .A(n31), .B(\CARRYB[10][6] ), .C(n32), .YC(\CARRYB[11][6] ), 
        .YS(\SUMB[11][6] ) );
  FAX1 S2_11_5 ( .A(n30), .B(\CARRYB[10][5] ), .C(\SUMB[10][6] ), .YC(
        \CARRYB[11][5] ), .YS(\SUMB[11][5] ) );
  FAX1 S3_10_6 ( .A(n31), .B(\CARRYB[9][6] ), .C(n32), .YC(\CARRYB[10][6] ), 
        .YS(\SUMB[10][6] ) );
  FAX1 S2_10_5 ( .A(n30), .B(\CARRYB[9][5] ), .C(\SUMB[9][6] ), .YC(
        \CARRYB[10][5] ), .YS(\SUMB[10][5] ) );
  FAX1 S3_9_6 ( .A(n31), .B(\CARRYB[8][6] ), .C(n32), .YC(\CARRYB[9][6] ), 
        .YS(\SUMB[9][6] ) );
  FAX1 S2_9_5 ( .A(n30), .B(\CARRYB[8][5] ), .C(\SUMB[8][6] ), .YC(
        \CARRYB[9][5] ), .YS(\SUMB[9][5] ) );
  FAX1 S3_8_6 ( .A(n31), .B(\CARRYB[7][6] ), .C(n32), .YC(\CARRYB[8][6] ), 
        .YS(\SUMB[8][6] ) );
  FAX1 S2_8_5 ( .A(n30), .B(\CARRYB[7][5] ), .C(\SUMB[7][6] ), .YC(
        \CARRYB[8][5] ), .YS(\SUMB[8][5] ) );
  FAX1 S3_7_6 ( .A(n31), .B(\CARRYB[6][6] ), .C(n32), .YC(\CARRYB[7][6] ), 
        .YS(\SUMB[7][6] ) );
  FAX1 S2_7_5 ( .A(n30), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S3_6_6 ( .A(n31), .B(\CARRYB[5][6] ), .C(n32), .YC(\CARRYB[6][6] ), 
        .YS(\SUMB[6][6] ) );
  FAX1 S2_6_5 ( .A(n30), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S3_5_6 ( .A(n31), .B(\CARRYB[4][6] ), .C(n32), .YC(\CARRYB[5][6] ), 
        .YS(\SUMB[5][6] ) );
  FAX1 S2_5_5 ( .A(n30), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S3_4_6 ( .A(n31), .B(\CARRYB[3][6] ), .C(n32), .YC(\CARRYB[4][6] ), 
        .YS(\SUMB[4][6] ) );
  FAX1 S2_4_5 ( .A(n30), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S3_3_6 ( .A(n31), .B(\CARRYB[2][6] ), .C(n32), .YC(\CARRYB[3][6] ), 
        .YS(\SUMB[3][6] ) );
  FAX1 S2_3_5 ( .A(n30), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S3_2_6 ( .A(n31), .B(n9), .C(n32), .YC(\CARRYB[2][6] ), .YS(
        \SUMB[2][6] ) );
  NAND2X1 U9 ( .A(B[7]), .B(A[9]), .Y(n10) );
  AND2X2 U8 ( .A(\ab[0][7] ), .B(n31), .Y(n9) );
  FAX1 S2_2_5 ( .A(n30), .B(n8), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), .YS(
        \SUMB[2][5] ) );
  XOR2X1 U25 ( .A(n31), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  NAND2X1 U11 ( .A(B[6]), .B(A[9]), .Y(n12) );
  AND2X2 U7 ( .A(\ab[0][6] ), .B(n30), .Y(n8) );
  NAND2X1 U13 ( .A(B[5]), .B(A[9]), .Y(n14) );
  INVX4 U10 ( .A(n10), .Y(n32) );
  INVX4 U12 ( .A(n12), .Y(n31) );
  INVX4 U14 ( .A(n14), .Y(n30) );
  INVX4 U16 ( .A(n16), .Y(n29) );
  INVX4 U18 ( .A(n18), .Y(n28) );
  INVX4 U20 ( .A(n20), .Y(n27) );
  INVX4 U22 ( .A(n22), .Y(n26) );
  INVX4 U24 ( .A(n24), .Y(n33) );
endmodule


module CannyEdge_DW02_mult_16 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n22), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n21), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n20), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n18), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n17), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n16), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n72), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n33), .B(\SUMB[3][1] ), .Y(n6) );
  AND2X2 U6 ( .A(n38), .B(\SUMB[3][2] ), .Y(n7) );
  AND2X2 U7 ( .A(n34), .B(\SUMB[3][3] ), .Y(n8) );
  AND2X2 U8 ( .A(n35), .B(\SUMB[3][4] ), .Y(n9) );
  AND2X2 U9 ( .A(n36), .B(\SUMB[3][5] ), .Y(n10) );
  AND2X2 U10 ( .A(n32), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n37), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n11), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[4][1] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n24), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n25), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n26), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n27), .B(\SUMB[5][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n39), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n33), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n38), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n34), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n35), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n36), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n37), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n6), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n7), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n8), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n9), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n10), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n39), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n24), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n32), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n75), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n74), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n71), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  NOR2X1 U114 ( .A(n81), .B(n80), .Y(\ab[2][7] ) );
  NOR2X1 U115 ( .A(n81), .B(n79), .Y(\ab[2][6] ) );
  NOR2X1 U116 ( .A(n81), .B(n78), .Y(\ab[2][5] ) );
  NOR2X1 U117 ( .A(n81), .B(n77), .Y(\ab[2][4] ) );
  NOR2X1 U118 ( .A(n81), .B(n76), .Y(\ab[2][3] ) );
  NOR2X1 U119 ( .A(n81), .B(n84), .Y(\ab[2][2] ) );
  NOR2X1 U120 ( .A(n81), .B(n73), .Y(\ab[2][1] ) );
  NOR2X1 U121 ( .A(n81), .B(n85), .Y(\ab[2][0] ) );
  NOR2X1 U122 ( .A(n80), .B(n82), .Y(\ab[1][7] ) );
  NOR2X1 U123 ( .A(n79), .B(n82), .Y(\ab[1][6] ) );
  NOR2X1 U124 ( .A(n78), .B(n82), .Y(\ab[1][5] ) );
  NOR2X1 U125 ( .A(n77), .B(n82), .Y(\ab[1][4] ) );
  NOR2X1 U126 ( .A(n76), .B(n82), .Y(\ab[1][3] ) );
  NOR2X1 U127 ( .A(n84), .B(n82), .Y(\ab[1][2] ) );
  NOR2X1 U128 ( .A(n73), .B(n82), .Y(\ab[1][1] ) );
  NOR2X1 U129 ( .A(n85), .B(n82), .Y(\ab[1][0] ) );
  NOR2X1 U130 ( .A(n80), .B(n83), .Y(\ab[0][7] ) );
  NOR2X1 U131 ( .A(n79), .B(n83), .Y(\ab[0][6] ) );
  NOR2X1 U132 ( .A(n78), .B(n83), .Y(\ab[0][5] ) );
  NOR2X1 U133 ( .A(n77), .B(n83), .Y(\ab[0][4] ) );
  NOR2X1 U134 ( .A(n76), .B(n83), .Y(\ab[0][3] ) );
  NOR2X1 U135 ( .A(n84), .B(n83), .Y(\ab[0][2] ) );
  NOR2X1 U136 ( .A(n73), .B(n83), .Y(\ab[0][1] ) );
  NOR2X1 U137 ( .A(n85), .B(n83), .Y(PRODUCT[0]) );
  INVX2 U99 ( .A(n49), .Y(n71) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n72) );
  INVX2 U101 ( .A(B[1]), .Y(n73) );
  INVX2 U102 ( .A(n52), .Y(n74) );
  INVX2 U103 ( .A(n48), .Y(n75) );
  INVX2 U104 ( .A(B[3]), .Y(n76) );
  INVX2 U105 ( .A(B[4]), .Y(n77) );
  INVX2 U106 ( .A(B[5]), .Y(n78) );
  INVX2 U107 ( .A(B[6]), .Y(n79) );
  INVX2 U108 ( .A(B[7]), .Y(n80) );
  INVX2 U109 ( .A(A[2]), .Y(n81) );
  INVX2 U110 ( .A(A[1]), .Y(n82) );
  INVX2 U111 ( .A(A[0]), .Y(n83) );
  INVX2 U112 ( .A(B[2]), .Y(n84) );
  INVX2 U113 ( .A(B[0]), .Y(n85) );
endmodule


module CannyEdge_DW01_add_39 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_17 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][7] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n61, n62, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n21), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n19), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n18), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n17), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n16), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n15), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(n23), .B(n67), .Y(n3) );
  AND2X2 U3 ( .A(n36), .B(\SUMB[3][2] ), .Y(n4) );
  AND2X2 U4 ( .A(n37), .B(\SUMB[3][3] ), .Y(n5) );
  AND2X2 U5 ( .A(n38), .B(\SUMB[3][4] ), .Y(n6) );
  AND2X2 U6 ( .A(n39), .B(\SUMB[3][5] ), .Y(n7) );
  AND2X2 U7 ( .A(n35), .B(\SUMB[6][1] ), .Y(n8) );
  AND2X2 U8 ( .A(n27), .B(\SUMB[6][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n28), .B(\SUMB[6][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n29), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n31), .B(\SUMB[6][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n40), .B(\CARRYB[2][6] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[4][1] ), .B(n34), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n13), .B(n67), .Y(n22) );
  AND2X2 U22 ( .A(n22), .B(n67), .Y(n23) );
  AND2X2 U23 ( .A(n4), .B(\SUMB[4][2] ), .Y(n24) );
  AND2X2 U24 ( .A(n5), .B(\SUMB[4][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n6), .B(\SUMB[4][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n24), .B(\SUMB[5][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n25), .B(\SUMB[5][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n26), .B(\SUMB[5][4] ), .Y(n29) );
  AND2X2 U29 ( .A(n7), .B(\SUMB[4][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n30), .B(\SUMB[5][5] ), .Y(n31) );
  AND2X2 U31 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[7][1] ), .B(n8), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[3][1] ), .B(n32), .Y(n34) );
  AND2X2 U34 ( .A(\SUMB[5][1] ), .B(n14), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n39) );
  AND2X2 U39 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n40) );
  AND2X2 U40 ( .A(QA), .B(QB), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n67), .Y(n42) );
  AND2X2 U42 ( .A(n67), .B(n3), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n9), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n11), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n12), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n8), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n9), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n10), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n12), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n67), .B(n3), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n41), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U55 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U56 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U57 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U58 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U59 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U60 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U61 ( .A(\SUMB[7][0] ), .B(n67), .Y(\A1[5] ) );
  XOR2X1 U62 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U63 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U64 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U65 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U66 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U67 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U68 ( .A(\SUMB[3][1] ), .B(n32), .Y(\A1[2] ) );
  XOR2X1 U69 ( .A(\SUMB[3][2] ), .B(n36), .Y(\SUMB[4][1] ) );
  XOR2X1 U70 ( .A(\SUMB[3][3] ), .B(n37), .Y(\SUMB[4][2] ) );
  XOR2X1 U71 ( .A(\SUMB[3][4] ), .B(n38), .Y(\SUMB[4][3] ) );
  XOR2X1 U72 ( .A(\SUMB[3][5] ), .B(n39), .Y(\SUMB[4][4] ) );
  XOR2X1 U73 ( .A(\CARRYB[2][6] ), .B(n40), .Y(\SUMB[4][5] ) );
  XOR2X1 U74 ( .A(\SUMB[4][1] ), .B(n34), .Y(\A1[3] ) );
  XOR2X1 U75 ( .A(\SUMB[4][2] ), .B(n4), .Y(\SUMB[5][1] ) );
  XOR2X1 U76 ( .A(\SUMB[4][3] ), .B(n5), .Y(\SUMB[5][2] ) );
  XOR2X1 U77 ( .A(\SUMB[4][4] ), .B(n6), .Y(\SUMB[5][3] ) );
  XOR2X1 U78 ( .A(\SUMB[4][5] ), .B(n7), .Y(\SUMB[5][4] ) );
  XOR2X1 U79 ( .A(n67), .B(n13), .Y(\SUMB[5][5] ) );
  XOR2X1 U80 ( .A(\SUMB[5][1] ), .B(n14), .Y(\A1[4] ) );
  XOR2X1 U81 ( .A(\SUMB[5][2] ), .B(n24), .Y(\SUMB[6][1] ) );
  XOR2X1 U82 ( .A(\SUMB[5][3] ), .B(n25), .Y(\SUMB[6][2] ) );
  XOR2X1 U83 ( .A(\SUMB[5][4] ), .B(n26), .Y(\SUMB[6][3] ) );
  XOR2X1 U84 ( .A(\SUMB[5][5] ), .B(n30), .Y(\SUMB[6][4] ) );
  XOR2X1 U85 ( .A(n67), .B(n22), .Y(\SUMB[6][5] ) );
  XOR2X1 U86 ( .A(\SUMB[6][1] ), .B(n35), .Y(\SUMB[7][0] ) );
  XOR2X1 U87 ( .A(\SUMB[6][2] ), .B(n27), .Y(\SUMB[7][1] ) );
  XOR2X1 U88 ( .A(\SUMB[6][3] ), .B(n28), .Y(\SUMB[7][2] ) );
  XOR2X1 U89 ( .A(\SUMB[6][4] ), .B(n29), .Y(\SUMB[7][3] ) );
  XOR2X1 U90 ( .A(\SUMB[6][5] ), .B(n31), .Y(\SUMB[7][4] ) );
  XOR2X1 U91 ( .A(n67), .B(n23), .Y(\SUMB[7][5] ) );
  XOR2X1 U92 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  NOR2X1 U105 ( .A(n66), .B(n73), .Y(\ab[2][6] ) );
  NOR2X1 U106 ( .A(n66), .B(n72), .Y(\ab[2][5] ) );
  NOR2X1 U107 ( .A(n66), .B(n71), .Y(\ab[2][4] ) );
  NOR2X1 U108 ( .A(n66), .B(n70), .Y(\ab[2][3] ) );
  NOR2X1 U109 ( .A(n66), .B(n69), .Y(\ab[2][2] ) );
  NOR2X1 U110 ( .A(n66), .B(n68), .Y(\ab[2][1] ) );
  NOR2X1 U111 ( .A(n66), .B(n75), .Y(\ab[2][0] ) );
  MUX2X1 U112 ( .B(n61), .A(n62), .S(A[1]), .Y(\ab[1][7] ) );
  NOR2X1 U113 ( .A(n73), .B(n76), .Y(\ab[1][6] ) );
  NOR2X1 U114 ( .A(n72), .B(n76), .Y(\ab[1][5] ) );
  NOR2X1 U115 ( .A(n71), .B(n76), .Y(\ab[1][4] ) );
  NOR2X1 U116 ( .A(n70), .B(n76), .Y(\ab[1][3] ) );
  NOR2X1 U117 ( .A(n69), .B(n76), .Y(\ab[1][2] ) );
  NOR2X1 U118 ( .A(n68), .B(n76), .Y(\ab[1][1] ) );
  NOR2X1 U119 ( .A(n75), .B(n76), .Y(\ab[1][0] ) );
  MUX2X1 U120 ( .B(n61), .A(n62), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U121 ( .A(B[7]), .B(n66), .Y(n62) );
  NOR2X1 U122 ( .A(n73), .B(n74), .Y(\ab[0][6] ) );
  NOR2X1 U123 ( .A(n72), .B(n74), .Y(\ab[0][5] ) );
  NOR2X1 U124 ( .A(n71), .B(n74), .Y(\ab[0][4] ) );
  NOR2X1 U125 ( .A(n70), .B(n74), .Y(\ab[0][3] ) );
  NOR2X1 U126 ( .A(n69), .B(n74), .Y(\ab[0][2] ) );
  NOR2X1 U127 ( .A(n68), .B(n74), .Y(\ab[0][1] ) );
  NAND2X1 U128 ( .A(QA), .B(B[7]), .Y(n61) );
  NOR2X1 U129 ( .A(B[7]), .B(n66), .Y(QB) );
  NOR2X1 U130 ( .A(n75), .B(n74), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_39 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n33, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n66) );
  INVX2 U97 ( .A(n61), .Y(n67) );
  INVX2 U98 ( .A(B[1]), .Y(n68) );
  INVX2 U99 ( .A(B[2]), .Y(n69) );
  INVX2 U100 ( .A(B[3]), .Y(n70) );
  INVX2 U101 ( .A(B[4]), .Y(n71) );
  INVX2 U102 ( .A(B[5]), .Y(n72) );
  INVX2 U103 ( .A(B[6]), .Y(n73) );
  INVX2 U104 ( .A(A[0]), .Y(n74) );
  INVX2 U131 ( .A(B[0]), .Y(n75) );
  INVX2 U132 ( .A(A[1]), .Y(n76) );
endmodule


module CannyEdge_DW01_add_40 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_18 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][7] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n61, n62, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n21), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n19), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n18), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n17), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n16), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n15), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(n23), .B(n67), .Y(n3) );
  AND2X2 U3 ( .A(n37), .B(\SUMB[3][2] ), .Y(n4) );
  AND2X2 U4 ( .A(n38), .B(\SUMB[3][3] ), .Y(n5) );
  AND2X2 U5 ( .A(n40), .B(\SUMB[3][4] ), .Y(n6) );
  AND2X2 U6 ( .A(n39), .B(\SUMB[3][5] ), .Y(n7) );
  AND2X2 U7 ( .A(n36), .B(\SUMB[6][1] ), .Y(n8) );
  AND2X2 U8 ( .A(n28), .B(\SUMB[6][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n29), .B(\SUMB[6][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n30), .B(\SUMB[6][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n32), .B(\SUMB[6][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n41), .B(\CARRYB[2][6] ), .Y(n13) );
  AND2X2 U13 ( .A(\SUMB[4][1] ), .B(n35), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n21) );
  AND2X2 U21 ( .A(n13), .B(n67), .Y(n22) );
  AND2X2 U22 ( .A(n22), .B(n67), .Y(n23) );
  AND2X2 U23 ( .A(QA), .B(QB), .Y(n24) );
  AND2X2 U24 ( .A(n4), .B(\SUMB[4][2] ), .Y(n25) );
  AND2X2 U25 ( .A(n5), .B(\SUMB[4][3] ), .Y(n26) );
  AND2X2 U26 ( .A(n6), .B(\SUMB[4][4] ), .Y(n27) );
  AND2X2 U27 ( .A(n25), .B(\SUMB[5][2] ), .Y(n28) );
  AND2X2 U28 ( .A(n26), .B(\SUMB[5][3] ), .Y(n29) );
  AND2X2 U29 ( .A(n27), .B(\SUMB[5][4] ), .Y(n30) );
  AND2X2 U30 ( .A(n7), .B(\SUMB[4][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n31), .B(\SUMB[5][5] ), .Y(n32) );
  AND2X2 U32 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n33) );
  AND2X2 U33 ( .A(\SUMB[7][1] ), .B(n8), .Y(n34) );
  AND2X2 U34 ( .A(\SUMB[3][1] ), .B(n33), .Y(n35) );
  AND2X2 U35 ( .A(\SUMB[5][1] ), .B(n14), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n39) );
  AND2X2 U39 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n40) );
  AND2X2 U40 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n67), .Y(n42) );
  AND2X2 U42 ( .A(n67), .B(n3), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n9), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n11), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n12), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n8), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n9), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n10), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n11), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n12), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n67), .B(n3), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n24), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U55 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U56 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U57 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U58 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U59 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U60 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U61 ( .A(\SUMB[7][0] ), .B(n67), .Y(\A1[5] ) );
  XOR2X1 U62 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U63 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U64 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U65 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U66 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U67 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U68 ( .A(\SUMB[3][1] ), .B(n33), .Y(\A1[2] ) );
  XOR2X1 U69 ( .A(\SUMB[3][2] ), .B(n37), .Y(\SUMB[4][1] ) );
  XOR2X1 U70 ( .A(\SUMB[3][3] ), .B(n38), .Y(\SUMB[4][2] ) );
  XOR2X1 U71 ( .A(\SUMB[3][4] ), .B(n40), .Y(\SUMB[4][3] ) );
  XOR2X1 U72 ( .A(\SUMB[3][5] ), .B(n39), .Y(\SUMB[4][4] ) );
  XOR2X1 U73 ( .A(\CARRYB[2][6] ), .B(n41), .Y(\SUMB[4][5] ) );
  XOR2X1 U74 ( .A(\SUMB[4][1] ), .B(n35), .Y(\A1[3] ) );
  XOR2X1 U75 ( .A(\SUMB[4][2] ), .B(n4), .Y(\SUMB[5][1] ) );
  XOR2X1 U76 ( .A(\SUMB[4][3] ), .B(n5), .Y(\SUMB[5][2] ) );
  XOR2X1 U77 ( .A(\SUMB[4][4] ), .B(n6), .Y(\SUMB[5][3] ) );
  XOR2X1 U78 ( .A(\SUMB[4][5] ), .B(n7), .Y(\SUMB[5][4] ) );
  XOR2X1 U79 ( .A(n67), .B(n13), .Y(\SUMB[5][5] ) );
  XOR2X1 U80 ( .A(\SUMB[5][1] ), .B(n14), .Y(\A1[4] ) );
  XOR2X1 U81 ( .A(\SUMB[5][2] ), .B(n25), .Y(\SUMB[6][1] ) );
  XOR2X1 U82 ( .A(\SUMB[5][3] ), .B(n26), .Y(\SUMB[6][2] ) );
  XOR2X1 U83 ( .A(\SUMB[5][4] ), .B(n27), .Y(\SUMB[6][3] ) );
  XOR2X1 U84 ( .A(\SUMB[5][5] ), .B(n31), .Y(\SUMB[6][4] ) );
  XOR2X1 U85 ( .A(n67), .B(n22), .Y(\SUMB[6][5] ) );
  XOR2X1 U86 ( .A(\SUMB[6][1] ), .B(n36), .Y(\SUMB[7][0] ) );
  XOR2X1 U87 ( .A(\SUMB[6][2] ), .B(n28), .Y(\SUMB[7][1] ) );
  XOR2X1 U88 ( .A(\SUMB[6][3] ), .B(n29), .Y(\SUMB[7][2] ) );
  XOR2X1 U89 ( .A(\SUMB[6][4] ), .B(n30), .Y(\SUMB[7][3] ) );
  XOR2X1 U90 ( .A(\SUMB[6][5] ), .B(n32), .Y(\SUMB[7][4] ) );
  XOR2X1 U91 ( .A(n67), .B(n23), .Y(\SUMB[7][5] ) );
  XOR2X1 U92 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  NOR2X1 U105 ( .A(n66), .B(n73), .Y(\ab[2][6] ) );
  NOR2X1 U106 ( .A(n66), .B(n72), .Y(\ab[2][5] ) );
  NOR2X1 U107 ( .A(n66), .B(n71), .Y(\ab[2][4] ) );
  NOR2X1 U108 ( .A(n66), .B(n70), .Y(\ab[2][3] ) );
  NOR2X1 U109 ( .A(n66), .B(n69), .Y(\ab[2][2] ) );
  NOR2X1 U110 ( .A(n66), .B(n68), .Y(\ab[2][1] ) );
  NOR2X1 U111 ( .A(n66), .B(n75), .Y(\ab[2][0] ) );
  MUX2X1 U112 ( .B(n61), .A(n62), .S(A[1]), .Y(\ab[1][7] ) );
  NOR2X1 U113 ( .A(n73), .B(n76), .Y(\ab[1][6] ) );
  NOR2X1 U114 ( .A(n72), .B(n76), .Y(\ab[1][5] ) );
  NOR2X1 U115 ( .A(n71), .B(n76), .Y(\ab[1][4] ) );
  NOR2X1 U116 ( .A(n70), .B(n76), .Y(\ab[1][3] ) );
  NOR2X1 U117 ( .A(n69), .B(n76), .Y(\ab[1][2] ) );
  NOR2X1 U118 ( .A(n68), .B(n76), .Y(\ab[1][1] ) );
  NOR2X1 U119 ( .A(n75), .B(n76), .Y(\ab[1][0] ) );
  MUX2X1 U120 ( .B(n61), .A(n62), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U121 ( .A(B[7]), .B(n66), .Y(n62) );
  NOR2X1 U122 ( .A(n73), .B(n74), .Y(\ab[0][6] ) );
  NOR2X1 U123 ( .A(n72), .B(n74), .Y(\ab[0][5] ) );
  NOR2X1 U124 ( .A(n71), .B(n74), .Y(\ab[0][4] ) );
  NOR2X1 U125 ( .A(n70), .B(n74), .Y(\ab[0][3] ) );
  NOR2X1 U126 ( .A(n69), .B(n74), .Y(\ab[0][2] ) );
  NOR2X1 U127 ( .A(n68), .B(n74), .Y(\ab[0][1] ) );
  NAND2X1 U128 ( .A(QA), .B(B[7]), .Y(n61) );
  NOR2X1 U129 ( .A(B[7]), .B(n66), .Y(QB) );
  NOR2X1 U130 ( .A(n75), .B(n74), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_40 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n34, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n66) );
  INVX2 U97 ( .A(n61), .Y(n67) );
  INVX2 U98 ( .A(B[1]), .Y(n68) );
  INVX2 U99 ( .A(B[2]), .Y(n69) );
  INVX2 U100 ( .A(B[3]), .Y(n70) );
  INVX2 U101 ( .A(B[4]), .Y(n71) );
  INVX2 U102 ( .A(B[5]), .Y(n72) );
  INVX2 U103 ( .A(B[6]), .Y(n73) );
  INVX2 U104 ( .A(A[0]), .Y(n74) );
  INVX2 U131 ( .A(B[0]), .Y(n75) );
  INVX2 U132 ( .A(A[1]), .Y(n76) );
endmodule


module CannyEdge_DW01_cmp2_3 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174;

  AND2X2 U1 ( .A(n130), .B(n60), .Y(n1) );
  MUX2X1 U59 ( .B(n1), .A(TC), .S(A[31]), .Y(GE_GT) );
  AOI21X1 U60 ( .A(A[29]), .B(n173), .C(n61), .Y(n60) );
  AOI21X1 U61 ( .A(B[29]), .B(n131), .C(n62), .Y(n61) );
  OAI21X1 U62 ( .A(A[28]), .B(n172), .C(n63), .Y(n62) );
  OAI21X1 U63 ( .A(B[28]), .B(n132), .C(n64), .Y(n63) );
  AOI21X1 U64 ( .A(A[27]), .B(n171), .C(n65), .Y(n64) );
  AOI21X1 U65 ( .A(B[27]), .B(n133), .C(n66), .Y(n65) );
  OAI21X1 U66 ( .A(A[26]), .B(n170), .C(n67), .Y(n66) );
  OAI21X1 U67 ( .A(B[26]), .B(n134), .C(n68), .Y(n67) );
  AOI21X1 U68 ( .A(A[25]), .B(n169), .C(n69), .Y(n68) );
  AOI21X1 U69 ( .A(B[25]), .B(n135), .C(n70), .Y(n69) );
  OAI21X1 U70 ( .A(A[24]), .B(n168), .C(n71), .Y(n70) );
  OAI21X1 U71 ( .A(B[24]), .B(n136), .C(n72), .Y(n71) );
  AOI21X1 U72 ( .A(A[23]), .B(n167), .C(n73), .Y(n72) );
  AOI21X1 U73 ( .A(B[23]), .B(n137), .C(n74), .Y(n73) );
  OAI21X1 U74 ( .A(A[22]), .B(n166), .C(n75), .Y(n74) );
  OAI21X1 U75 ( .A(B[22]), .B(n138), .C(n76), .Y(n75) );
  AOI21X1 U76 ( .A(A[21]), .B(n165), .C(n77), .Y(n76) );
  AOI21X1 U77 ( .A(B[21]), .B(n139), .C(n78), .Y(n77) );
  OAI21X1 U78 ( .A(A[20]), .B(n164), .C(n79), .Y(n78) );
  OAI21X1 U79 ( .A(B[20]), .B(n140), .C(n80), .Y(n79) );
  AOI21X1 U80 ( .A(A[19]), .B(n163), .C(n81), .Y(n80) );
  AOI21X1 U81 ( .A(B[19]), .B(n141), .C(n82), .Y(n81) );
  OAI21X1 U82 ( .A(A[18]), .B(n162), .C(n83), .Y(n82) );
  OAI21X1 U83 ( .A(B[18]), .B(n142), .C(n84), .Y(n83) );
  AOI21X1 U84 ( .A(A[17]), .B(n161), .C(n85), .Y(n84) );
  AOI21X1 U85 ( .A(B[17]), .B(n143), .C(n86), .Y(n85) );
  OAI21X1 U86 ( .A(A[16]), .B(n160), .C(n87), .Y(n86) );
  OAI21X1 U87 ( .A(B[16]), .B(n144), .C(n88), .Y(n87) );
  AOI21X1 U88 ( .A(A[15]), .B(n159), .C(n89), .Y(n88) );
  AOI21X1 U89 ( .A(B[15]), .B(n145), .C(n90), .Y(n89) );
  OAI21X1 U90 ( .A(A[14]), .B(n158), .C(n91), .Y(n90) );
  OAI21X1 U91 ( .A(B[14]), .B(n146), .C(n92), .Y(n91) );
  AOI21X1 U92 ( .A(A[13]), .B(n157), .C(n93), .Y(n92) );
  AOI21X1 U93 ( .A(B[13]), .B(n147), .C(n94), .Y(n93) );
  OAI21X1 U94 ( .A(A[12]), .B(n156), .C(n95), .Y(n94) );
  OAI21X1 U95 ( .A(B[12]), .B(n148), .C(n96), .Y(n95) );
  AOI21X1 U96 ( .A(A[11]), .B(n155), .C(n97), .Y(n96) );
  AOI21X1 U97 ( .A(B[11]), .B(n149), .C(n98), .Y(n97) );
  OAI21X1 U98 ( .A(A[10]), .B(n154), .C(n99), .Y(n98) );
  OAI21X1 U99 ( .A(B[9]), .B(n128), .C(n100), .Y(n99) );
  AOI21X1 U100 ( .A(A[10]), .B(n154), .C(n101), .Y(n100) );
  AOI21X1 U101 ( .A(B[9]), .B(n128), .C(n102), .Y(n101) );
  OAI21X1 U102 ( .A(A[8]), .B(n174), .C(n103), .Y(n102) );
  OAI21X1 U103 ( .A(B[8]), .B(n129), .C(n104), .Y(n103) );
  AOI21X1 U104 ( .A(A[7]), .B(n118), .C(n105), .Y(n104) );
  AOI21X1 U105 ( .A(B[7]), .B(n150), .C(n106), .Y(n105) );
  OAI21X1 U106 ( .A(A[6]), .B(n119), .C(n107), .Y(n106) );
  OAI21X1 U107 ( .A(B[6]), .B(n151), .C(n108), .Y(n107) );
  AOI21X1 U108 ( .A(A[5]), .B(n120), .C(n109), .Y(n108) );
  AOI21X1 U109 ( .A(B[5]), .B(n152), .C(n110), .Y(n109) );
  OAI21X1 U110 ( .A(A[4]), .B(n121), .C(n111), .Y(n110) );
  OAI21X1 U111 ( .A(B[4]), .B(n153), .C(n112), .Y(n111) );
  AOI21X1 U112 ( .A(A[3]), .B(n122), .C(n113), .Y(n112) );
  AOI21X1 U113 ( .A(B[3]), .B(n127), .C(n114), .Y(n113) );
  OAI21X1 U114 ( .A(A[2]), .B(n123), .C(n115), .Y(n114) );
  OAI21X1 U115 ( .A(B[2]), .B(n126), .C(n116), .Y(n115) );
  AOI22X1 U116 ( .A(n117), .B(A[0]), .C(A[1]), .D(n124), .Y(n116) );
  AOI21X1 U117 ( .A(B[1]), .B(n125), .C(B[0]), .Y(n117) );
  INVX2 U2 ( .A(B[7]), .Y(n118) );
  INVX2 U3 ( .A(B[6]), .Y(n119) );
  INVX2 U4 ( .A(B[5]), .Y(n120) );
  INVX2 U5 ( .A(B[4]), .Y(n121) );
  INVX2 U6 ( .A(B[3]), .Y(n122) );
  INVX2 U7 ( .A(B[2]), .Y(n123) );
  INVX2 U8 ( .A(B[1]), .Y(n124) );
  INVX2 U9 ( .A(A[1]), .Y(n125) );
  INVX2 U10 ( .A(A[2]), .Y(n126) );
  INVX2 U11 ( .A(A[3]), .Y(n127) );
  INVX2 U12 ( .A(A[9]), .Y(n128) );
  INVX2 U13 ( .A(A[8]), .Y(n129) );
  INVX2 U14 ( .A(A[30]), .Y(n130) );
  INVX2 U15 ( .A(A[29]), .Y(n131) );
  INVX2 U16 ( .A(A[28]), .Y(n132) );
  INVX2 U17 ( .A(A[27]), .Y(n133) );
  INVX2 U18 ( .A(A[26]), .Y(n134) );
  INVX2 U19 ( .A(A[25]), .Y(n135) );
  INVX2 U20 ( .A(A[24]), .Y(n136) );
  INVX2 U21 ( .A(A[23]), .Y(n137) );
  INVX2 U22 ( .A(A[22]), .Y(n138) );
  INVX2 U23 ( .A(A[21]), .Y(n139) );
  INVX2 U24 ( .A(A[20]), .Y(n140) );
  INVX2 U25 ( .A(A[19]), .Y(n141) );
  INVX2 U26 ( .A(A[18]), .Y(n142) );
  INVX2 U27 ( .A(A[17]), .Y(n143) );
  INVX2 U28 ( .A(A[16]), .Y(n144) );
  INVX2 U29 ( .A(A[15]), .Y(n145) );
  INVX2 U30 ( .A(A[14]), .Y(n146) );
  INVX2 U31 ( .A(A[13]), .Y(n147) );
  INVX2 U32 ( .A(A[12]), .Y(n148) );
  INVX2 U33 ( .A(A[11]), .Y(n149) );
  INVX2 U34 ( .A(A[7]), .Y(n150) );
  INVX2 U35 ( .A(A[6]), .Y(n151) );
  INVX2 U36 ( .A(A[5]), .Y(n152) );
  INVX2 U37 ( .A(A[4]), .Y(n153) );
  INVX2 U38 ( .A(B[10]), .Y(n154) );
  INVX2 U39 ( .A(B[11]), .Y(n155) );
  INVX2 U40 ( .A(B[12]), .Y(n156) );
  INVX2 U41 ( .A(B[13]), .Y(n157) );
  INVX2 U42 ( .A(B[14]), .Y(n158) );
  INVX2 U43 ( .A(B[15]), .Y(n159) );
  INVX2 U44 ( .A(B[16]), .Y(n160) );
  INVX2 U45 ( .A(B[17]), .Y(n161) );
  INVX2 U46 ( .A(B[18]), .Y(n162) );
  INVX2 U47 ( .A(B[19]), .Y(n163) );
  INVX2 U48 ( .A(B[20]), .Y(n164) );
  INVX2 U49 ( .A(B[21]), .Y(n165) );
  INVX2 U50 ( .A(B[22]), .Y(n166) );
  INVX2 U51 ( .A(B[23]), .Y(n167) );
  INVX2 U52 ( .A(B[24]), .Y(n168) );
  INVX2 U53 ( .A(B[25]), .Y(n169) );
  INVX2 U54 ( .A(B[26]), .Y(n170) );
  INVX2 U55 ( .A(B[27]), .Y(n171) );
  INVX2 U56 ( .A(B[28]), .Y(n172) );
  INVX2 U57 ( .A(B[29]), .Y(n173) );
  INVX2 U58 ( .A(B[8]), .Y(n174) );
endmodule


module CannyEdge_DW01_add_41 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n141, n142, n143, n144, n145, n146, n147,
         n148, n149;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U31 ( .A(n30), .B(n31), .Y(SUM[9]) );
  NOR2X1 U32 ( .A(n130), .B(n32), .Y(n31) );
  XOR2X1 U33 ( .A(n34), .B(n134), .Y(SUM[8]) );
  NAND2X1 U34 ( .A(n133), .B(n35), .Y(n34) );
  XOR2X1 U35 ( .A(n37), .B(n38), .Y(SUM[7]) );
  XOR2X1 U36 ( .A(n135), .B(B[7]), .Y(n38) );
  OAI21X1 U37 ( .A(B[6]), .B(A[6]), .C(n37), .Y(n39) );
  XOR2X1 U38 ( .A(n40), .B(n41), .Y(SUM[29]) );
  XOR2X1 U39 ( .A(B[29]), .B(A[29]), .Y(n41) );
  OAI21X1 U40 ( .A(n42), .B(n43), .C(n44), .Y(n40) );
  XOR2X1 U41 ( .A(n45), .B(n43), .Y(SUM[28]) );
  AOI21X1 U42 ( .A(n137), .B(n46), .C(n47), .Y(n43) );
  NAND2X1 U43 ( .A(n136), .B(n44), .Y(n45) );
  NAND2X1 U44 ( .A(B[28]), .B(A[28]), .Y(n44) );
  NOR2X1 U45 ( .A(B[28]), .B(A[28]), .Y(n42) );
  XOR2X1 U46 ( .A(n46), .B(n49), .Y(SUM[27]) );
  NOR2X1 U47 ( .A(n47), .B(n48), .Y(n49) );
  NOR2X1 U48 ( .A(B[27]), .B(A[27]), .Y(n48) );
  AND2X1 U49 ( .A(B[27]), .B(A[27]), .Y(n47) );
  OAI21X1 U50 ( .A(n50), .B(n51), .C(n52), .Y(n46) );
  XOR2X1 U51 ( .A(n53), .B(n51), .Y(SUM[26]) );
  AOI21X1 U52 ( .A(n139), .B(n54), .C(n55), .Y(n51) );
  NAND2X1 U53 ( .A(n138), .B(n52), .Y(n53) );
  NAND2X1 U54 ( .A(B[26]), .B(A[26]), .Y(n52) );
  NOR2X1 U55 ( .A(B[26]), .B(A[26]), .Y(n50) );
  XOR2X1 U56 ( .A(n54), .B(n57), .Y(SUM[25]) );
  NOR2X1 U57 ( .A(n55), .B(n56), .Y(n57) );
  NOR2X1 U58 ( .A(B[25]), .B(A[25]), .Y(n56) );
  AND2X1 U59 ( .A(B[25]), .B(A[25]), .Y(n55) );
  OAI21X1 U60 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  XOR2X1 U61 ( .A(n61), .B(n59), .Y(SUM[24]) );
  AOI21X1 U62 ( .A(n143), .B(n62), .C(n63), .Y(n59) );
  NAND2X1 U63 ( .A(n142), .B(n60), .Y(n61) );
  NAND2X1 U64 ( .A(B[24]), .B(A[24]), .Y(n60) );
  NOR2X1 U65 ( .A(B[24]), .B(A[24]), .Y(n58) );
  XOR2X1 U66 ( .A(n62), .B(n65), .Y(SUM[23]) );
  NOR2X1 U67 ( .A(n63), .B(n64), .Y(n65) );
  NOR2X1 U68 ( .A(B[23]), .B(A[23]), .Y(n64) );
  AND2X1 U69 ( .A(B[23]), .B(A[23]), .Y(n63) );
  OAI21X1 U70 ( .A(n66), .B(n67), .C(n68), .Y(n62) );
  XOR2X1 U71 ( .A(n69), .B(n67), .Y(SUM[22]) );
  AOI21X1 U72 ( .A(n145), .B(n70), .C(n71), .Y(n67) );
  NAND2X1 U73 ( .A(n144), .B(n68), .Y(n69) );
  NAND2X1 U74 ( .A(B[22]), .B(A[22]), .Y(n68) );
  NOR2X1 U75 ( .A(B[22]), .B(A[22]), .Y(n66) );
  XOR2X1 U76 ( .A(n70), .B(n73), .Y(SUM[21]) );
  NOR2X1 U77 ( .A(n71), .B(n72), .Y(n73) );
  NOR2X1 U78 ( .A(B[21]), .B(A[21]), .Y(n72) );
  AND2X1 U79 ( .A(B[21]), .B(A[21]), .Y(n71) );
  OAI21X1 U80 ( .A(n74), .B(n75), .C(n76), .Y(n70) );
  XOR2X1 U81 ( .A(n77), .B(n75), .Y(SUM[20]) );
  AOI21X1 U82 ( .A(n147), .B(n78), .C(n79), .Y(n75) );
  NAND2X1 U83 ( .A(n146), .B(n76), .Y(n77) );
  NAND2X1 U84 ( .A(B[20]), .B(A[20]), .Y(n76) );
  NOR2X1 U85 ( .A(B[20]), .B(A[20]), .Y(n74) );
  XOR2X1 U86 ( .A(n78), .B(n81), .Y(SUM[19]) );
  NOR2X1 U87 ( .A(n79), .B(n80), .Y(n81) );
  NOR2X1 U88 ( .A(B[19]), .B(A[19]), .Y(n80) );
  AND2X1 U89 ( .A(B[19]), .B(A[19]), .Y(n79) );
  OAI21X1 U90 ( .A(n82), .B(n83), .C(n84), .Y(n78) );
  XOR2X1 U91 ( .A(n85), .B(n83), .Y(SUM[18]) );
  AOI21X1 U92 ( .A(n149), .B(n86), .C(n87), .Y(n83) );
  NAND2X1 U93 ( .A(n148), .B(n84), .Y(n85) );
  NAND2X1 U94 ( .A(B[18]), .B(A[18]), .Y(n84) );
  NOR2X1 U95 ( .A(B[18]), .B(A[18]), .Y(n82) );
  XOR2X1 U96 ( .A(n86), .B(n89), .Y(SUM[17]) );
  NOR2X1 U97 ( .A(n87), .B(n88), .Y(n89) );
  NOR2X1 U98 ( .A(B[17]), .B(A[17]), .Y(n88) );
  AND2X1 U99 ( .A(B[17]), .B(A[17]), .Y(n87) );
  OAI21X1 U100 ( .A(n90), .B(n91), .C(n92), .Y(n86) );
  XOR2X1 U101 ( .A(n93), .B(n91), .Y(SUM[16]) );
  AOI21X1 U102 ( .A(n122), .B(n94), .C(n95), .Y(n91) );
  NAND2X1 U103 ( .A(n121), .B(n92), .Y(n93) );
  NAND2X1 U104 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NOR2X1 U105 ( .A(B[16]), .B(A[16]), .Y(n90) );
  XOR2X1 U106 ( .A(n94), .B(n97), .Y(SUM[15]) );
  NOR2X1 U107 ( .A(n95), .B(n96), .Y(n97) );
  NOR2X1 U108 ( .A(B[15]), .B(A[15]), .Y(n96) );
  AND2X1 U109 ( .A(B[15]), .B(A[15]), .Y(n95) );
  OAI21X1 U110 ( .A(n98), .B(n99), .C(n100), .Y(n94) );
  XOR2X1 U111 ( .A(n101), .B(n99), .Y(SUM[14]) );
  AOI21X1 U112 ( .A(n124), .B(n102), .C(n103), .Y(n99) );
  NAND2X1 U113 ( .A(n123), .B(n100), .Y(n101) );
  NAND2X1 U114 ( .A(B[14]), .B(A[14]), .Y(n100) );
  NOR2X1 U115 ( .A(B[14]), .B(A[14]), .Y(n98) );
  XOR2X1 U116 ( .A(n102), .B(n105), .Y(SUM[13]) );
  NOR2X1 U117 ( .A(n103), .B(n104), .Y(n105) );
  NOR2X1 U118 ( .A(B[13]), .B(A[13]), .Y(n104) );
  AND2X1 U119 ( .A(B[13]), .B(A[13]), .Y(n103) );
  OAI21X1 U120 ( .A(n106), .B(n126), .C(n107), .Y(n102) );
  XOR2X1 U121 ( .A(n108), .B(n126), .Y(SUM[12]) );
  OAI21X1 U122 ( .A(n110), .B(n111), .C(n112), .Y(n109) );
  AOI21X1 U123 ( .A(n113), .B(n129), .C(n128), .Y(n111) );
  NAND2X1 U124 ( .A(n125), .B(n107), .Y(n108) );
  NAND2X1 U125 ( .A(B[12]), .B(A[12]), .Y(n107) );
  NOR2X1 U126 ( .A(B[12]), .B(A[12]), .Y(n106) );
  XOR2X1 U127 ( .A(n115), .B(n116), .Y(SUM[11]) );
  NOR2X1 U128 ( .A(n127), .B(n110), .Y(n116) );
  NOR2X1 U129 ( .A(B[11]), .B(A[11]), .Y(n110) );
  NAND2X1 U130 ( .A(B[11]), .B(A[11]), .Y(n112) );
  OAI21X1 U131 ( .A(n117), .B(n131), .C(n114), .Y(n115) );
  XOR2X1 U132 ( .A(n118), .B(n131), .Y(SUM[10]) );
  OAI21X1 U133 ( .A(n132), .B(n32), .C(n33), .Y(n113) );
  NAND2X1 U134 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NOR2X1 U135 ( .A(B[9]), .B(A[9]), .Y(n32) );
  OAI21X1 U136 ( .A(n36), .B(n134), .C(n35), .Y(n30) );
  NAND2X1 U137 ( .A(B[8]), .B(A[8]), .Y(n35) );
  OAI21X1 U138 ( .A(n37), .B(n135), .C(n120), .Y(n119) );
  OAI21X1 U139 ( .A(n141), .B(A[7]), .C(B[7]), .Y(n120) );
  NAND2X1 U140 ( .A(B[6]), .B(A[6]), .Y(n37) );
  NOR2X1 U141 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NAND2X1 U142 ( .A(n129), .B(n114), .Y(n118) );
  NAND2X1 U143 ( .A(B[10]), .B(A[10]), .Y(n114) );
  NOR2X1 U144 ( .A(B[10]), .B(A[10]), .Y(n117) );
  INVX2 U2 ( .A(n90), .Y(n121) );
  INVX2 U3 ( .A(n96), .Y(n122) );
  INVX2 U4 ( .A(n98), .Y(n123) );
  INVX2 U5 ( .A(n104), .Y(n124) );
  INVX2 U6 ( .A(n106), .Y(n125) );
  INVX2 U7 ( .A(n109), .Y(n126) );
  INVX2 U8 ( .A(n112), .Y(n127) );
  INVX2 U9 ( .A(n114), .Y(n128) );
  INVX2 U10 ( .A(n117), .Y(n129) );
  INVX2 U11 ( .A(n33), .Y(n130) );
  INVX2 U12 ( .A(n113), .Y(n131) );
  INVX2 U13 ( .A(n30), .Y(n132) );
  INVX2 U14 ( .A(n36), .Y(n133) );
  INVX2 U15 ( .A(n119), .Y(n134) );
  INVX2 U16 ( .A(A[7]), .Y(n135) );
  INVX2 U17 ( .A(n42), .Y(n136) );
  INVX2 U18 ( .A(n48), .Y(n137) );
  INVX2 U19 ( .A(n50), .Y(n138) );
  INVX2 U20 ( .A(n56), .Y(n139) );
  INVX2 U21 ( .A(n39), .Y(SUM[6]) );
  INVX2 U22 ( .A(n37), .Y(n141) );
  INVX2 U23 ( .A(n58), .Y(n142) );
  INVX2 U24 ( .A(n64), .Y(n143) );
  INVX2 U25 ( .A(n66), .Y(n144) );
  INVX2 U26 ( .A(n72), .Y(n145) );
  INVX2 U27 ( .A(n74), .Y(n146) );
  INVX2 U28 ( .A(n80), .Y(n147) );
  INVX2 U29 ( .A(n82), .Y(n148) );
  INVX2 U30 ( .A(n88), .Y(n149) );
endmodule


module CannyEdge_DW02_mult_19 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] , \ab[7][27] ,
         \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][31] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][31] , \ab[3][30] ,
         \ab[3][29] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] , \ab[2][27] ,
         \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][31] ,
         \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] ,
         \ab[0][25] , \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] ,
         \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] ,
         \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] ,
         \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] ,
         \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] ,
         \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[30] , n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n110, n111, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S14_31_0 ( .A(n117), .B(\CARRYB[7][23] ), .C(\SUMB[7][24] ), .YC(
        \A2[30] ), .YS(\A1[29] ) );
  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S4_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S4_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S4_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S4_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  FAX1 S4_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S4_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S4_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S4_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  FAX1 S4_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S4_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S4_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S4_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  FAX1 S4_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S4_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S4_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S4_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  FAX1 S4_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S4_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S4_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S4_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  FAX1 S4_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S4_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S5_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .C(\ab[6][31] ), .YC(
        \CARRYB[7][30] ), .YS(\SUMB[7][30] ) );
  FAX1 S14_31 ( .A(QA), .B(QB), .C(\ab[7][31] ), .YC(\CARRYB[7][31] ), .YS(
        \SUMB[7][31] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  FAX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  FAX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  FAX1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  FAX1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  FAX1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .C(\ab[5][31] ), .YC(
        \CARRYB[6][30] ), .YS(\SUMB[6][30] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .C(\ab[4][31] ), .YC(
        \CARRYB[5][30] ), .YS(\SUMB[5][30] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .C(\ab[3][31] ), .YC(
        \CARRYB[4][30] ), .YS(\SUMB[4][30] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .C(\ab[2][31] ), .YC(
        \CARRYB[3][30] ), .YS(\SUMB[3][30] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n42), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n41), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n40), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n39), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n38), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n37), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n36), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n35), .C(\SUMB[1][8] ), .YC(\CARRYB[2][7] ), 
        .YS(\SUMB[2][7] ) );
  FAX1 S2_2_8 ( .A(\ab[2][8] ), .B(n34), .C(\SUMB[1][9] ), .YC(\CARRYB[2][8] ), 
        .YS(\SUMB[2][8] ) );
  FAX1 S2_2_9 ( .A(\ab[2][9] ), .B(n33), .C(\SUMB[1][10] ), .YC(\CARRYB[2][9] ), .YS(\SUMB[2][9] ) );
  FAX1 S2_2_10 ( .A(\ab[2][10] ), .B(n32), .C(\SUMB[1][11] ), .YC(
        \CARRYB[2][10] ), .YS(\SUMB[2][10] ) );
  FAX1 S2_2_11 ( .A(\ab[2][11] ), .B(n31), .C(\SUMB[1][12] ), .YC(
        \CARRYB[2][11] ), .YS(\SUMB[2][11] ) );
  FAX1 S2_2_12 ( .A(\ab[2][12] ), .B(n30), .C(\SUMB[1][13] ), .YC(
        \CARRYB[2][12] ), .YS(\SUMB[2][12] ) );
  FAX1 S2_2_13 ( .A(\ab[2][13] ), .B(n29), .C(\SUMB[1][14] ), .YC(
        \CARRYB[2][13] ), .YS(\SUMB[2][13] ) );
  FAX1 S2_2_14 ( .A(\ab[2][14] ), .B(n28), .C(\SUMB[1][15] ), .YC(
        \CARRYB[2][14] ), .YS(\SUMB[2][14] ) );
  FAX1 S2_2_15 ( .A(\ab[2][15] ), .B(n27), .C(\SUMB[1][16] ), .YC(
        \CARRYB[2][15] ), .YS(\SUMB[2][15] ) );
  FAX1 S2_2_16 ( .A(\ab[2][16] ), .B(n26), .C(\SUMB[1][17] ), .YC(
        \CARRYB[2][16] ), .YS(\SUMB[2][16] ) );
  FAX1 S2_2_17 ( .A(\ab[2][17] ), .B(n25), .C(\SUMB[1][18] ), .YC(
        \CARRYB[2][17] ), .YS(\SUMB[2][17] ) );
  FAX1 S2_2_18 ( .A(\ab[2][18] ), .B(n24), .C(\SUMB[1][19] ), .YC(
        \CARRYB[2][18] ), .YS(\SUMB[2][18] ) );
  FAX1 S2_2_19 ( .A(\ab[2][19] ), .B(n23), .C(\SUMB[1][20] ), .YC(
        \CARRYB[2][19] ), .YS(\SUMB[2][19] ) );
  FAX1 S2_2_20 ( .A(\ab[2][20] ), .B(n22), .C(\SUMB[1][21] ), .YC(
        \CARRYB[2][20] ), .YS(\SUMB[2][20] ) );
  FAX1 S2_2_21 ( .A(\ab[2][21] ), .B(n21), .C(\SUMB[1][22] ), .YC(
        \CARRYB[2][21] ), .YS(\SUMB[2][21] ) );
  FAX1 S2_2_22 ( .A(\ab[2][22] ), .B(n20), .C(\SUMB[1][23] ), .YC(
        \CARRYB[2][22] ), .YS(\SUMB[2][22] ) );
  FAX1 S2_2_23 ( .A(\ab[2][23] ), .B(n19), .C(\SUMB[1][24] ), .YC(
        \CARRYB[2][23] ), .YS(\SUMB[2][23] ) );
  FAX1 S2_2_24 ( .A(\ab[2][24] ), .B(n18), .C(\SUMB[1][25] ), .YC(
        \CARRYB[2][24] ), .YS(\SUMB[2][24] ) );
  FAX1 S2_2_25 ( .A(\ab[2][25] ), .B(n17), .C(\SUMB[1][26] ), .YC(
        \CARRYB[2][25] ), .YS(\SUMB[2][25] ) );
  FAX1 S2_2_26 ( .A(\ab[2][26] ), .B(n16), .C(\SUMB[1][27] ), .YC(
        \CARRYB[2][26] ), .YS(\SUMB[2][26] ) );
  FAX1 S2_2_27 ( .A(\ab[2][27] ), .B(n15), .C(\SUMB[1][28] ), .YC(
        \CARRYB[2][27] ), .YS(\SUMB[2][27] ) );
  FAX1 S2_2_28 ( .A(\ab[2][28] ), .B(n14), .C(\SUMB[1][29] ), .YC(
        \CARRYB[2][28] ), .YS(\SUMB[2][28] ) );
  FAX1 S2_2_29 ( .A(\ab[2][29] ), .B(n13), .C(\SUMB[1][30] ), .YC(
        \CARRYB[2][29] ), .YS(\SUMB[2][29] ) );
  FAX1 S3_2_30 ( .A(\ab[2][30] ), .B(n12), .C(\ab[1][31] ), .YC(
        \CARRYB[2][30] ), .YS(\SUMB[2][30] ) );
  AND2X2 U2 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(n3) );
  AND2X2 U3 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(n4) );
  AND2X2 U4 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(n5) );
  AND2X2 U5 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(n6) );
  AND2X2 U6 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(n7) );
  AND2X2 U7 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(n8) );
  AND2X2 U8 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(n9) );
  AND2X2 U9 ( .A(TC), .B(A[7]), .Y(n10) );
  AND2X2 U10 ( .A(A[7]), .B(n115), .Y(n11) );
  AND2X2 U11 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Y(n12) );
  AND2X2 U12 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Y(n13) );
  AND2X2 U13 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Y(n24) );
  AND2X2 U24 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Y(n25) );
  AND2X2 U25 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Y(n26) );
  AND2X2 U26 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Y(n27) );
  AND2X2 U27 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n28) );
  AND2X2 U28 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n29) );
  AND2X2 U29 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n30) );
  AND2X2 U30 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Y(n31) );
  AND2X2 U31 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n36) );
  AND2X2 U36 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n37) );
  AND2X2 U37 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n38) );
  AND2X2 U38 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n39) );
  AND2X2 U39 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n40) );
  AND2X2 U40 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n41) );
  AND2X2 U41 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n42) );
  AND2X2 U42 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][0] ), .B(n10), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(n53) );
  AND2X2 U53 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(n54) );
  AND2X2 U54 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(n55) );
  AND2X2 U55 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(n56) );
  AND2X2 U56 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(n57) );
  AND2X2 U57 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(n58) );
  AND2X2 U58 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(n59) );
  AND2X2 U59 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(n60) );
  AND2X2 U60 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(n61) );
  AND2X2 U61 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(n62) );
  AND2X2 U62 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(n63) );
  AND2X2 U63 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n64) );
  AND2X2 U64 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(n65) );
  AND2X2 U65 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(n66) );
  XOR2X1 U68 ( .A(\SUMB[7][0] ), .B(n10), .Y(\A1[5] ) );
  XOR2X1 U69 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  XOR2X1 U70 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  XOR2X1 U71 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  XOR2X1 U72 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  XOR2X1 U73 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  XOR2X1 U74 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  XOR2X1 U75 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  XOR2X1 U76 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  XOR2X1 U77 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  XOR2X1 U78 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  XOR2X1 U79 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  XOR2X1 U80 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  XOR2X1 U81 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  XOR2X1 U82 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  XOR2X1 U83 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  XOR2X1 U84 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  XOR2X1 U85 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  XOR2X1 U86 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  XOR2X1 U87 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  XOR2X1 U88 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  XOR2X1 U89 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  XOR2X1 U90 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  XOR2X1 U91 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  XOR2X1 U92 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  XOR2X1 U93 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  XOR2X1 U94 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  XOR2X1 U95 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  XOR2X1 U96 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  XOR2X1 U97 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  XOR2X1 U98 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(\A1[36] ) );
  XOR2X1 U99 ( .A(\CARRYB[7][31] ), .B(TC), .Y(\A1[37] ) );
  XOR2X1 U100 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U101 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U102 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U103 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U104 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U105 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U106 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U107 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  XOR2X1 U108 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(\SUMB[1][8] ) );
  XOR2X1 U109 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Y(\SUMB[1][9] ) );
  XOR2X1 U110 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Y(\SUMB[1][10] ) );
  XOR2X1 U111 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U112 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Y(\SUMB[1][12] ) );
  XOR2X1 U113 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  XOR2X1 U114 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  XOR2X1 U115 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Y(\SUMB[1][15] ) );
  XOR2X1 U116 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Y(\SUMB[1][16] ) );
  XOR2X1 U117 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Y(\SUMB[1][17] ) );
  XOR2X1 U118 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Y(\SUMB[1][18] ) );
  XOR2X1 U119 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Y(\SUMB[1][19] ) );
  XOR2X1 U120 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Y(\SUMB[1][20] ) );
  XOR2X1 U121 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Y(\SUMB[1][21] ) );
  XOR2X1 U122 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Y(\SUMB[1][22] ) );
  XOR2X1 U123 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Y(\SUMB[1][23] ) );
  XOR2X1 U124 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Y(\SUMB[1][24] ) );
  XOR2X1 U125 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Y(\SUMB[1][25] ) );
  XOR2X1 U126 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Y(\SUMB[1][26] ) );
  XOR2X1 U127 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Y(\SUMB[1][27] ) );
  XOR2X1 U128 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Y(\SUMB[1][28] ) );
  XOR2X1 U129 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Y(\SUMB[1][29] ) );
  XOR2X1 U130 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Y(\SUMB[1][30] ) );
  MUX2X1 U171 ( .B(n116), .A(n114), .S(B[9]), .Y(\ab[7][9] ) );
  MUX2X1 U172 ( .B(n116), .A(n114), .S(B[8]), .Y(\ab[7][8] ) );
  MUX2X1 U173 ( .B(n116), .A(n114), .S(B[7]), .Y(\ab[7][7] ) );
  MUX2X1 U174 ( .B(n116), .A(n114), .S(B[6]), .Y(\ab[7][6] ) );
  MUX2X1 U175 ( .B(n116), .A(n114), .S(B[5]), .Y(\ab[7][5] ) );
  MUX2X1 U176 ( .B(n116), .A(n114), .S(B[4]), .Y(\ab[7][4] ) );
  MUX2X1 U177 ( .B(n116), .A(n114), .S(B[3]), .Y(\ab[7][3] ) );
  AND2X1 U178 ( .A(A[7]), .B(B[31]), .Y(\ab[7][31] ) );
  MUX2X1 U179 ( .B(n116), .A(n114), .S(B[30]), .Y(\ab[7][30] ) );
  MUX2X1 U180 ( .B(n116), .A(n114), .S(B[2]), .Y(\ab[7][2] ) );
  MUX2X1 U181 ( .B(n116), .A(n114), .S(B[29]), .Y(\ab[7][29] ) );
  MUX2X1 U182 ( .B(n116), .A(n114), .S(B[28]), .Y(\ab[7][28] ) );
  MUX2X1 U183 ( .B(n116), .A(n114), .S(B[27]), .Y(\ab[7][27] ) );
  MUX2X1 U184 ( .B(n116), .A(n114), .S(B[26]), .Y(\ab[7][26] ) );
  MUX2X1 U185 ( .B(n116), .A(n114), .S(B[25]), .Y(\ab[7][25] ) );
  MUX2X1 U186 ( .B(n116), .A(n114), .S(B[24]), .Y(\ab[7][24] ) );
  MUX2X1 U187 ( .B(n116), .A(n114), .S(B[23]), .Y(\ab[7][23] ) );
  MUX2X1 U188 ( .B(n116), .A(n114), .S(B[22]), .Y(\ab[7][22] ) );
  MUX2X1 U189 ( .B(n116), .A(n114), .S(B[21]), .Y(\ab[7][21] ) );
  MUX2X1 U190 ( .B(n116), .A(n114), .S(B[20]), .Y(\ab[7][20] ) );
  MUX2X1 U191 ( .B(n116), .A(n114), .S(B[1]), .Y(\ab[7][1] ) );
  MUX2X1 U192 ( .B(n116), .A(n114), .S(B[19]), .Y(\ab[7][19] ) );
  MUX2X1 U193 ( .B(n116), .A(n114), .S(B[18]), .Y(\ab[7][18] ) );
  MUX2X1 U194 ( .B(n116), .A(n114), .S(B[17]), .Y(\ab[7][17] ) );
  MUX2X1 U195 ( .B(n116), .A(n114), .S(B[16]), .Y(\ab[7][16] ) );
  MUX2X1 U196 ( .B(n116), .A(n114), .S(B[15]), .Y(\ab[7][15] ) );
  MUX2X1 U197 ( .B(n116), .A(n114), .S(B[14]), .Y(\ab[7][14] ) );
  MUX2X1 U198 ( .B(n116), .A(n114), .S(B[13]), .Y(\ab[7][13] ) );
  MUX2X1 U199 ( .B(n116), .A(n114), .S(B[12]), .Y(\ab[7][12] ) );
  MUX2X1 U200 ( .B(n116), .A(n114), .S(B[11]), .Y(\ab[7][11] ) );
  MUX2X1 U201 ( .B(n116), .A(n114), .S(B[10]), .Y(\ab[7][10] ) );
  MUX2X1 U202 ( .B(n116), .A(n114), .S(B[0]), .Y(\ab[7][0] ) );
  NOR2X1 U203 ( .A(n154), .B(n123), .Y(\ab[6][9] ) );
  NOR2X1 U204 ( .A(n153), .B(n123), .Y(\ab[6][8] ) );
  NOR2X1 U205 ( .A(n152), .B(n123), .Y(\ab[6][7] ) );
  NOR2X1 U206 ( .A(n151), .B(n123), .Y(\ab[6][6] ) );
  NOR2X1 U207 ( .A(n150), .B(n123), .Y(\ab[6][5] ) );
  NOR2X1 U208 ( .A(n149), .B(n123), .Y(\ab[6][4] ) );
  NOR2X1 U209 ( .A(n147), .B(n123), .Y(\ab[6][3] ) );
  MUX2X1 U210 ( .B(n110), .A(n111), .S(A[6]), .Y(\ab[6][31] ) );
  NOR2X1 U211 ( .A(n148), .B(n123), .Y(\ab[6][30] ) );
  NOR2X1 U212 ( .A(n136), .B(n123), .Y(\ab[6][2] ) );
  NOR2X1 U213 ( .A(n146), .B(n123), .Y(\ab[6][29] ) );
  NOR2X1 U214 ( .A(n145), .B(n123), .Y(\ab[6][28] ) );
  NOR2X1 U215 ( .A(n144), .B(n123), .Y(\ab[6][27] ) );
  NOR2X1 U216 ( .A(n143), .B(n123), .Y(\ab[6][26] ) );
  NOR2X1 U217 ( .A(n142), .B(n123), .Y(\ab[6][25] ) );
  NOR2X1 U218 ( .A(n141), .B(n123), .Y(\ab[6][24] ) );
  NOR2X1 U219 ( .A(n140), .B(n123), .Y(\ab[6][23] ) );
  NOR2X1 U220 ( .A(n139), .B(n123), .Y(\ab[6][22] ) );
  NOR2X1 U221 ( .A(n138), .B(n123), .Y(\ab[6][21] ) );
  NOR2X1 U222 ( .A(n137), .B(n123), .Y(\ab[6][20] ) );
  NOR2X1 U223 ( .A(n125), .B(n123), .Y(\ab[6][1] ) );
  NOR2X1 U224 ( .A(n135), .B(n123), .Y(\ab[6][19] ) );
  NOR2X1 U225 ( .A(n134), .B(n123), .Y(\ab[6][18] ) );
  NOR2X1 U226 ( .A(n133), .B(n123), .Y(\ab[6][17] ) );
  NOR2X1 U227 ( .A(n132), .B(n123), .Y(\ab[6][16] ) );
  NOR2X1 U228 ( .A(n131), .B(n123), .Y(\ab[6][15] ) );
  NOR2X1 U229 ( .A(n130), .B(n123), .Y(\ab[6][14] ) );
  NOR2X1 U230 ( .A(n129), .B(n123), .Y(\ab[6][13] ) );
  NOR2X1 U231 ( .A(n128), .B(n123), .Y(\ab[6][12] ) );
  NOR2X1 U232 ( .A(n127), .B(n123), .Y(\ab[6][11] ) );
  NOR2X1 U233 ( .A(n126), .B(n123), .Y(\ab[6][10] ) );
  NOR2X1 U234 ( .A(n124), .B(n123), .Y(\ab[6][0] ) );
  NOR2X1 U235 ( .A(n154), .B(n122), .Y(\ab[5][9] ) );
  NOR2X1 U236 ( .A(n153), .B(n122), .Y(\ab[5][8] ) );
  NOR2X1 U237 ( .A(n152), .B(n122), .Y(\ab[5][7] ) );
  NOR2X1 U238 ( .A(n151), .B(n122), .Y(\ab[5][6] ) );
  NOR2X1 U239 ( .A(n150), .B(n122), .Y(\ab[5][5] ) );
  NOR2X1 U240 ( .A(n149), .B(n122), .Y(\ab[5][4] ) );
  NOR2X1 U241 ( .A(n147), .B(n122), .Y(\ab[5][3] ) );
  MUX2X1 U242 ( .B(n110), .A(n111), .S(A[5]), .Y(\ab[5][31] ) );
  NOR2X1 U243 ( .A(n148), .B(n122), .Y(\ab[5][30] ) );
  NOR2X1 U244 ( .A(n136), .B(n122), .Y(\ab[5][2] ) );
  NOR2X1 U245 ( .A(n146), .B(n122), .Y(\ab[5][29] ) );
  NOR2X1 U246 ( .A(n145), .B(n122), .Y(\ab[5][28] ) );
  NOR2X1 U247 ( .A(n144), .B(n122), .Y(\ab[5][27] ) );
  NOR2X1 U248 ( .A(n143), .B(n122), .Y(\ab[5][26] ) );
  NOR2X1 U249 ( .A(n142), .B(n122), .Y(\ab[5][25] ) );
  NOR2X1 U250 ( .A(n141), .B(n122), .Y(\ab[5][24] ) );
  NOR2X1 U251 ( .A(n140), .B(n122), .Y(\ab[5][23] ) );
  NOR2X1 U252 ( .A(n139), .B(n122), .Y(\ab[5][22] ) );
  NOR2X1 U253 ( .A(n138), .B(n122), .Y(\ab[5][21] ) );
  NOR2X1 U254 ( .A(n137), .B(n122), .Y(\ab[5][20] ) );
  NOR2X1 U255 ( .A(n125), .B(n122), .Y(\ab[5][1] ) );
  NOR2X1 U256 ( .A(n135), .B(n122), .Y(\ab[5][19] ) );
  NOR2X1 U257 ( .A(n134), .B(n122), .Y(\ab[5][18] ) );
  NOR2X1 U258 ( .A(n133), .B(n122), .Y(\ab[5][17] ) );
  NOR2X1 U259 ( .A(n132), .B(n122), .Y(\ab[5][16] ) );
  NOR2X1 U260 ( .A(n131), .B(n122), .Y(\ab[5][15] ) );
  NOR2X1 U261 ( .A(n130), .B(n122), .Y(\ab[5][14] ) );
  NOR2X1 U262 ( .A(n129), .B(n122), .Y(\ab[5][13] ) );
  NOR2X1 U263 ( .A(n128), .B(n122), .Y(\ab[5][12] ) );
  NOR2X1 U264 ( .A(n127), .B(n122), .Y(\ab[5][11] ) );
  NOR2X1 U265 ( .A(n126), .B(n122), .Y(\ab[5][10] ) );
  NOR2X1 U266 ( .A(n124), .B(n122), .Y(\ab[5][0] ) );
  NOR2X1 U267 ( .A(n154), .B(n121), .Y(\ab[4][9] ) );
  NOR2X1 U268 ( .A(n153), .B(n121), .Y(\ab[4][8] ) );
  NOR2X1 U269 ( .A(n152), .B(n121), .Y(\ab[4][7] ) );
  NOR2X1 U270 ( .A(n151), .B(n121), .Y(\ab[4][6] ) );
  NOR2X1 U271 ( .A(n150), .B(n121), .Y(\ab[4][5] ) );
  NOR2X1 U272 ( .A(n149), .B(n121), .Y(\ab[4][4] ) );
  NOR2X1 U273 ( .A(n147), .B(n121), .Y(\ab[4][3] ) );
  MUX2X1 U274 ( .B(n110), .A(n111), .S(A[4]), .Y(\ab[4][31] ) );
  NOR2X1 U275 ( .A(n148), .B(n121), .Y(\ab[4][30] ) );
  NOR2X1 U276 ( .A(n136), .B(n121), .Y(\ab[4][2] ) );
  NOR2X1 U277 ( .A(n146), .B(n121), .Y(\ab[4][29] ) );
  NOR2X1 U278 ( .A(n145), .B(n121), .Y(\ab[4][28] ) );
  NOR2X1 U279 ( .A(n144), .B(n121), .Y(\ab[4][27] ) );
  NOR2X1 U280 ( .A(n143), .B(n121), .Y(\ab[4][26] ) );
  NOR2X1 U281 ( .A(n142), .B(n121), .Y(\ab[4][25] ) );
  NOR2X1 U282 ( .A(n141), .B(n121), .Y(\ab[4][24] ) );
  NOR2X1 U283 ( .A(n140), .B(n121), .Y(\ab[4][23] ) );
  NOR2X1 U284 ( .A(n139), .B(n121), .Y(\ab[4][22] ) );
  NOR2X1 U285 ( .A(n138), .B(n121), .Y(\ab[4][21] ) );
  NOR2X1 U286 ( .A(n137), .B(n121), .Y(\ab[4][20] ) );
  NOR2X1 U287 ( .A(n125), .B(n121), .Y(\ab[4][1] ) );
  NOR2X1 U288 ( .A(n135), .B(n121), .Y(\ab[4][19] ) );
  NOR2X1 U289 ( .A(n134), .B(n121), .Y(\ab[4][18] ) );
  NOR2X1 U290 ( .A(n133), .B(n121), .Y(\ab[4][17] ) );
  NOR2X1 U291 ( .A(n132), .B(n121), .Y(\ab[4][16] ) );
  NOR2X1 U292 ( .A(n131), .B(n121), .Y(\ab[4][15] ) );
  NOR2X1 U293 ( .A(n130), .B(n121), .Y(\ab[4][14] ) );
  NOR2X1 U294 ( .A(n129), .B(n121), .Y(\ab[4][13] ) );
  NOR2X1 U295 ( .A(n128), .B(n121), .Y(\ab[4][12] ) );
  NOR2X1 U296 ( .A(n127), .B(n121), .Y(\ab[4][11] ) );
  NOR2X1 U297 ( .A(n126), .B(n121), .Y(\ab[4][10] ) );
  NOR2X1 U298 ( .A(n124), .B(n121), .Y(\ab[4][0] ) );
  NOR2X1 U299 ( .A(n154), .B(n120), .Y(\ab[3][9] ) );
  NOR2X1 U300 ( .A(n153), .B(n120), .Y(\ab[3][8] ) );
  NOR2X1 U301 ( .A(n152), .B(n120), .Y(\ab[3][7] ) );
  NOR2X1 U302 ( .A(n151), .B(n120), .Y(\ab[3][6] ) );
  NOR2X1 U303 ( .A(n150), .B(n120), .Y(\ab[3][5] ) );
  NOR2X1 U304 ( .A(n149), .B(n120), .Y(\ab[3][4] ) );
  NOR2X1 U305 ( .A(n147), .B(n120), .Y(\ab[3][3] ) );
  MUX2X1 U306 ( .B(n110), .A(n111), .S(A[3]), .Y(\ab[3][31] ) );
  NOR2X1 U307 ( .A(n148), .B(n120), .Y(\ab[3][30] ) );
  NOR2X1 U308 ( .A(n136), .B(n120), .Y(\ab[3][2] ) );
  NOR2X1 U309 ( .A(n146), .B(n120), .Y(\ab[3][29] ) );
  NOR2X1 U310 ( .A(n145), .B(n120), .Y(\ab[3][28] ) );
  NOR2X1 U311 ( .A(n144), .B(n120), .Y(\ab[3][27] ) );
  NOR2X1 U312 ( .A(n143), .B(n120), .Y(\ab[3][26] ) );
  NOR2X1 U313 ( .A(n142), .B(n120), .Y(\ab[3][25] ) );
  NOR2X1 U314 ( .A(n141), .B(n120), .Y(\ab[3][24] ) );
  NOR2X1 U315 ( .A(n140), .B(n120), .Y(\ab[3][23] ) );
  NOR2X1 U316 ( .A(n139), .B(n120), .Y(\ab[3][22] ) );
  NOR2X1 U317 ( .A(n138), .B(n120), .Y(\ab[3][21] ) );
  NOR2X1 U318 ( .A(n137), .B(n120), .Y(\ab[3][20] ) );
  NOR2X1 U319 ( .A(n125), .B(n120), .Y(\ab[3][1] ) );
  NOR2X1 U320 ( .A(n135), .B(n120), .Y(\ab[3][19] ) );
  NOR2X1 U321 ( .A(n134), .B(n120), .Y(\ab[3][18] ) );
  NOR2X1 U322 ( .A(n133), .B(n120), .Y(\ab[3][17] ) );
  NOR2X1 U323 ( .A(n132), .B(n120), .Y(\ab[3][16] ) );
  NOR2X1 U324 ( .A(n131), .B(n120), .Y(\ab[3][15] ) );
  NOR2X1 U325 ( .A(n130), .B(n120), .Y(\ab[3][14] ) );
  NOR2X1 U326 ( .A(n129), .B(n120), .Y(\ab[3][13] ) );
  NOR2X1 U327 ( .A(n128), .B(n120), .Y(\ab[3][12] ) );
  NOR2X1 U328 ( .A(n127), .B(n120), .Y(\ab[3][11] ) );
  NOR2X1 U329 ( .A(n126), .B(n120), .Y(\ab[3][10] ) );
  NOR2X1 U330 ( .A(n124), .B(n120), .Y(\ab[3][0] ) );
  NOR2X1 U331 ( .A(n154), .B(n155), .Y(\ab[2][9] ) );
  NOR2X1 U332 ( .A(n153), .B(n155), .Y(\ab[2][8] ) );
  NOR2X1 U333 ( .A(n152), .B(n155), .Y(\ab[2][7] ) );
  NOR2X1 U334 ( .A(n151), .B(n155), .Y(\ab[2][6] ) );
  NOR2X1 U335 ( .A(n150), .B(n155), .Y(\ab[2][5] ) );
  NOR2X1 U336 ( .A(n149), .B(n155), .Y(\ab[2][4] ) );
  NOR2X1 U337 ( .A(n147), .B(n155), .Y(\ab[2][3] ) );
  MUX2X1 U338 ( .B(n110), .A(n111), .S(A[2]), .Y(\ab[2][31] ) );
  NOR2X1 U339 ( .A(n148), .B(n155), .Y(\ab[2][30] ) );
  NOR2X1 U340 ( .A(n136), .B(n155), .Y(\ab[2][2] ) );
  NOR2X1 U341 ( .A(n146), .B(n155), .Y(\ab[2][29] ) );
  NOR2X1 U342 ( .A(n145), .B(n155), .Y(\ab[2][28] ) );
  NOR2X1 U343 ( .A(n144), .B(n155), .Y(\ab[2][27] ) );
  NOR2X1 U344 ( .A(n143), .B(n155), .Y(\ab[2][26] ) );
  NOR2X1 U345 ( .A(n142), .B(n155), .Y(\ab[2][25] ) );
  NOR2X1 U346 ( .A(n141), .B(n155), .Y(\ab[2][24] ) );
  NOR2X1 U347 ( .A(n140), .B(n155), .Y(\ab[2][23] ) );
  NOR2X1 U348 ( .A(n139), .B(n155), .Y(\ab[2][22] ) );
  NOR2X1 U349 ( .A(n138), .B(n155), .Y(\ab[2][21] ) );
  NOR2X1 U350 ( .A(n137), .B(n155), .Y(\ab[2][20] ) );
  NOR2X1 U351 ( .A(n125), .B(n155), .Y(\ab[2][1] ) );
  NOR2X1 U352 ( .A(n135), .B(n155), .Y(\ab[2][19] ) );
  NOR2X1 U353 ( .A(n134), .B(n155), .Y(\ab[2][18] ) );
  NOR2X1 U354 ( .A(n133), .B(n155), .Y(\ab[2][17] ) );
  NOR2X1 U355 ( .A(n132), .B(n155), .Y(\ab[2][16] ) );
  NOR2X1 U356 ( .A(n131), .B(n155), .Y(\ab[2][15] ) );
  NOR2X1 U357 ( .A(n130), .B(n155), .Y(\ab[2][14] ) );
  NOR2X1 U358 ( .A(n129), .B(n155), .Y(\ab[2][13] ) );
  NOR2X1 U359 ( .A(n128), .B(n155), .Y(\ab[2][12] ) );
  NOR2X1 U360 ( .A(n127), .B(n155), .Y(\ab[2][11] ) );
  NOR2X1 U361 ( .A(n126), .B(n155), .Y(\ab[2][10] ) );
  NOR2X1 U362 ( .A(n124), .B(n155), .Y(\ab[2][0] ) );
  NOR2X1 U363 ( .A(n154), .B(n119), .Y(\ab[1][9] ) );
  NOR2X1 U364 ( .A(n153), .B(n119), .Y(\ab[1][8] ) );
  NOR2X1 U365 ( .A(n152), .B(n119), .Y(\ab[1][7] ) );
  NOR2X1 U366 ( .A(n151), .B(n119), .Y(\ab[1][6] ) );
  NOR2X1 U367 ( .A(n150), .B(n119), .Y(\ab[1][5] ) );
  NOR2X1 U368 ( .A(n149), .B(n119), .Y(\ab[1][4] ) );
  NOR2X1 U369 ( .A(n147), .B(n119), .Y(\ab[1][3] ) );
  MUX2X1 U370 ( .B(n110), .A(n111), .S(A[1]), .Y(\ab[1][31] ) );
  NOR2X1 U371 ( .A(n148), .B(n119), .Y(\ab[1][30] ) );
  NOR2X1 U372 ( .A(n136), .B(n119), .Y(\ab[1][2] ) );
  NOR2X1 U373 ( .A(n146), .B(n119), .Y(\ab[1][29] ) );
  NOR2X1 U374 ( .A(n145), .B(n119), .Y(\ab[1][28] ) );
  NOR2X1 U375 ( .A(n144), .B(n119), .Y(\ab[1][27] ) );
  NOR2X1 U376 ( .A(n143), .B(n119), .Y(\ab[1][26] ) );
  NOR2X1 U377 ( .A(n142), .B(n119), .Y(\ab[1][25] ) );
  NOR2X1 U378 ( .A(n141), .B(n119), .Y(\ab[1][24] ) );
  NOR2X1 U379 ( .A(n140), .B(n119), .Y(\ab[1][23] ) );
  NOR2X1 U380 ( .A(n139), .B(n119), .Y(\ab[1][22] ) );
  NOR2X1 U381 ( .A(n138), .B(n119), .Y(\ab[1][21] ) );
  NOR2X1 U382 ( .A(n137), .B(n119), .Y(\ab[1][20] ) );
  NOR2X1 U383 ( .A(n125), .B(n119), .Y(\ab[1][1] ) );
  NOR2X1 U384 ( .A(n135), .B(n119), .Y(\ab[1][19] ) );
  NOR2X1 U385 ( .A(n134), .B(n119), .Y(\ab[1][18] ) );
  NOR2X1 U386 ( .A(n133), .B(n119), .Y(\ab[1][17] ) );
  NOR2X1 U387 ( .A(n132), .B(n119), .Y(\ab[1][16] ) );
  NOR2X1 U388 ( .A(n131), .B(n119), .Y(\ab[1][15] ) );
  NOR2X1 U389 ( .A(n130), .B(n119), .Y(\ab[1][14] ) );
  NOR2X1 U390 ( .A(n129), .B(n119), .Y(\ab[1][13] ) );
  NOR2X1 U391 ( .A(n128), .B(n119), .Y(\ab[1][12] ) );
  NOR2X1 U392 ( .A(n127), .B(n119), .Y(\ab[1][11] ) );
  NOR2X1 U393 ( .A(n126), .B(n119), .Y(\ab[1][10] ) );
  NOR2X1 U394 ( .A(n124), .B(n119), .Y(\ab[1][0] ) );
  NOR2X1 U395 ( .A(n154), .B(n118), .Y(\ab[0][9] ) );
  NOR2X1 U396 ( .A(n153), .B(n118), .Y(\ab[0][8] ) );
  NOR2X1 U397 ( .A(n152), .B(n118), .Y(\ab[0][7] ) );
  NOR2X1 U398 ( .A(n151), .B(n118), .Y(\ab[0][6] ) );
  NOR2X1 U399 ( .A(n150), .B(n118), .Y(\ab[0][5] ) );
  NOR2X1 U400 ( .A(n149), .B(n118), .Y(\ab[0][4] ) );
  NOR2X1 U401 ( .A(n147), .B(n118), .Y(\ab[0][3] ) );
  MUX2X1 U402 ( .B(n110), .A(n111), .S(A[0]), .Y(\ab[0][31] ) );
  NAND2X1 U403 ( .A(B[31]), .B(n115), .Y(n111) );
  NOR2X1 U404 ( .A(n148), .B(n118), .Y(\ab[0][30] ) );
  NOR2X1 U405 ( .A(n136), .B(n118), .Y(\ab[0][2] ) );
  NOR2X1 U406 ( .A(n146), .B(n118), .Y(\ab[0][29] ) );
  NOR2X1 U407 ( .A(n145), .B(n118), .Y(\ab[0][28] ) );
  NOR2X1 U408 ( .A(n144), .B(n118), .Y(\ab[0][27] ) );
  NOR2X1 U409 ( .A(n143), .B(n118), .Y(\ab[0][26] ) );
  NOR2X1 U410 ( .A(n142), .B(n118), .Y(\ab[0][25] ) );
  NOR2X1 U411 ( .A(n141), .B(n118), .Y(\ab[0][24] ) );
  NOR2X1 U412 ( .A(n140), .B(n118), .Y(\ab[0][23] ) );
  NOR2X1 U413 ( .A(n139), .B(n118), .Y(\ab[0][22] ) );
  NOR2X1 U414 ( .A(n138), .B(n118), .Y(\ab[0][21] ) );
  NOR2X1 U415 ( .A(n137), .B(n118), .Y(\ab[0][20] ) );
  NOR2X1 U416 ( .A(n125), .B(n118), .Y(\ab[0][1] ) );
  NOR2X1 U417 ( .A(n135), .B(n118), .Y(\ab[0][19] ) );
  NOR2X1 U418 ( .A(n134), .B(n118), .Y(\ab[0][18] ) );
  NOR2X1 U419 ( .A(n133), .B(n118), .Y(\ab[0][17] ) );
  NOR2X1 U420 ( .A(n132), .B(n118), .Y(\ab[0][16] ) );
  NOR2X1 U421 ( .A(n131), .B(n118), .Y(\ab[0][15] ) );
  NOR2X1 U422 ( .A(n130), .B(n118), .Y(\ab[0][14] ) );
  NOR2X1 U423 ( .A(n129), .B(n118), .Y(\ab[0][13] ) );
  NOR2X1 U424 ( .A(n128), .B(n118), .Y(\ab[0][12] ) );
  NOR2X1 U425 ( .A(n127), .B(n118), .Y(\ab[0][11] ) );
  NOR2X1 U426 ( .A(n126), .B(n118), .Y(\ab[0][10] ) );
  NAND2X1 U427 ( .A(B[31]), .B(TC), .Y(n110) );
  NOR2X1 U428 ( .A(B[31]), .B(n115), .Y(QB) );
  NOR2X1 U429 ( .A(A[7]), .B(n115), .Y(QA) );
  NOR2X1 U430 ( .A(n124), .B(n118), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_41 FS_1 ( .A({\A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n9, n8, n7, 
        n6, n5, n4, n3, \A2[30] , n45, n54, n46, n55, n47, n56, n48, n57, n49, 
        n58, n50, n59, n51, n60, n52, n61, n53, n62, n63, n66, n64, n65, n43, 
        n44, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  INVX2 U131 ( .A(n11), .Y(n114) );
  INVX2 U132 ( .A(TC), .Y(n115) );
  INVX2 U133 ( .A(n10), .Y(n116) );
  INVX2 U134 ( .A(n110), .Y(n117) );
  INVX2 U135 ( .A(A[0]), .Y(n118) );
  INVX2 U136 ( .A(A[1]), .Y(n119) );
  INVX2 U137 ( .A(A[3]), .Y(n120) );
  INVX2 U138 ( .A(A[4]), .Y(n121) );
  INVX2 U139 ( .A(A[5]), .Y(n122) );
  INVX2 U140 ( .A(A[6]), .Y(n123) );
  INVX2 U141 ( .A(B[0]), .Y(n124) );
  INVX2 U142 ( .A(B[1]), .Y(n125) );
  INVX2 U143 ( .A(B[10]), .Y(n126) );
  INVX2 U144 ( .A(B[11]), .Y(n127) );
  INVX2 U145 ( .A(B[12]), .Y(n128) );
  INVX2 U146 ( .A(B[13]), .Y(n129) );
  INVX2 U147 ( .A(B[14]), .Y(n130) );
  INVX2 U148 ( .A(B[15]), .Y(n131) );
  INVX2 U149 ( .A(B[16]), .Y(n132) );
  INVX2 U150 ( .A(B[17]), .Y(n133) );
  INVX2 U151 ( .A(B[18]), .Y(n134) );
  INVX2 U152 ( .A(B[19]), .Y(n135) );
  INVX2 U153 ( .A(B[2]), .Y(n136) );
  INVX2 U154 ( .A(B[20]), .Y(n137) );
  INVX2 U155 ( .A(B[21]), .Y(n138) );
  INVX2 U156 ( .A(B[22]), .Y(n139) );
  INVX2 U157 ( .A(B[23]), .Y(n140) );
  INVX2 U158 ( .A(B[24]), .Y(n141) );
  INVX2 U159 ( .A(B[25]), .Y(n142) );
  INVX2 U160 ( .A(B[26]), .Y(n143) );
  INVX2 U161 ( .A(B[27]), .Y(n144) );
  INVX2 U162 ( .A(B[28]), .Y(n145) );
  INVX2 U163 ( .A(B[29]), .Y(n146) );
  INVX2 U164 ( .A(B[3]), .Y(n147) );
  INVX2 U165 ( .A(B[30]), .Y(n148) );
  INVX2 U166 ( .A(B[4]), .Y(n149) );
  INVX2 U167 ( .A(B[5]), .Y(n150) );
  INVX2 U168 ( .A(B[6]), .Y(n151) );
  INVX2 U169 ( .A(B[7]), .Y(n152) );
  INVX2 U170 ( .A(B[8]), .Y(n153) );
  INVX2 U431 ( .A(B[9]), .Y(n154) );
  INVX2 U432 ( .A(A[2]), .Y(n155) );
endmodule


module CannyEdge_DW01_cmp2_4 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188;

  MUX2X1 U63 ( .B(n63), .A(n64), .S(B[31]), .Y(GE_GT) );
  MUX2X1 U64 ( .B(TC), .A(n65), .S(A[31]), .Y(n64) );
  NOR2X1 U65 ( .A(n66), .B(n167), .Y(n65) );
  MUX2X1 U66 ( .B(n67), .A(n188), .S(A[31]), .Y(n63) );
  NAND2X1 U67 ( .A(n66), .B(n167), .Y(n67) );
  OAI21X1 U68 ( .A(A[29]), .B(n147), .C(n68), .Y(n66) );
  OAI21X1 U69 ( .A(B[29]), .B(n168), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(A[28]), .B(n146), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(B[28]), .B(n169), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(A[27]), .B(n145), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(B[27]), .B(n170), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(A[26]), .B(n144), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(B[26]), .B(n171), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(A[25]), .B(n143), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(B[25]), .B(n172), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(A[24]), .B(n142), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(B[24]), .B(n173), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(A[23]), .B(n141), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(B[23]), .B(n174), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(A[22]), .B(n140), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(B[22]), .B(n175), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(A[21]), .B(n139), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(B[21]), .B(n176), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(A[20]), .B(n138), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(B[20]), .B(n177), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(A[19]), .B(n137), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(B[19]), .B(n178), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(A[18]), .B(n136), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(B[18]), .B(n179), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(A[17]), .B(n135), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(B[17]), .B(n180), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(A[16]), .B(n148), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(B[16]), .B(n181), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(A[15]), .B(n149), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(B[15]), .B(n182), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(A[14]), .B(n150), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(B[14]), .B(n183), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(A[13]), .B(n151), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(B[13]), .B(n184), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(A[12]), .B(n152), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(B[12]), .B(n185), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(A[11]), .B(n153), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(B[11]), .B(n186), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(A[10]), .B(n154), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(B[10]), .B(n187), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(A[9]), .B(n155), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(B[9]), .B(n165), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(A[8]), .B(n156), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(B[8]), .B(n166), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(A[7]), .B(n157), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(B[7]), .B(n134), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(A[6]), .B(n158), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(B[6]), .B(n133), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(A[5]), .B(n159), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(B[5]), .B(n132), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(A[4]), .B(n160), .C(n118), .Y(n117) );
  AOI21X1 U119 ( .A(B[4]), .B(n131), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(A[3]), .B(n161), .C(n120), .Y(n119) );
  OAI21X1 U121 ( .A(B[3]), .B(n130), .C(n121), .Y(n120) );
  AOI21X1 U122 ( .A(A[2]), .B(n162), .C(n122), .Y(n121) );
  AOI21X1 U123 ( .A(B[2]), .B(n129), .C(n123), .Y(n122) );
  OAI21X1 U124 ( .A(A[1]), .B(n163), .C(n124), .Y(n123) );
  OAI21X1 U125 ( .A(B[1]), .B(n128), .C(n125), .Y(n124) );
  AOI21X1 U126 ( .A(A[0]), .B(n164), .C(n126), .Y(n125) );
  AOI21X1 U127 ( .A(B[0]), .B(n127), .C(LEQ), .Y(n126) );
  INVX2 U1 ( .A(A[0]), .Y(n127) );
  INVX2 U2 ( .A(A[1]), .Y(n128) );
  INVX2 U3 ( .A(A[2]), .Y(n129) );
  INVX2 U4 ( .A(A[3]), .Y(n130) );
  INVX2 U5 ( .A(A[4]), .Y(n131) );
  INVX2 U6 ( .A(A[5]), .Y(n132) );
  INVX2 U7 ( .A(A[6]), .Y(n133) );
  INVX2 U8 ( .A(A[7]), .Y(n134) );
  INVX2 U9 ( .A(B[17]), .Y(n135) );
  INVX2 U10 ( .A(B[18]), .Y(n136) );
  INVX2 U11 ( .A(B[19]), .Y(n137) );
  INVX2 U12 ( .A(B[20]), .Y(n138) );
  INVX2 U13 ( .A(B[21]), .Y(n139) );
  INVX2 U14 ( .A(B[22]), .Y(n140) );
  INVX2 U15 ( .A(B[23]), .Y(n141) );
  INVX2 U16 ( .A(B[24]), .Y(n142) );
  INVX2 U17 ( .A(B[25]), .Y(n143) );
  INVX2 U18 ( .A(B[26]), .Y(n144) );
  INVX2 U19 ( .A(B[27]), .Y(n145) );
  INVX2 U20 ( .A(B[28]), .Y(n146) );
  INVX2 U21 ( .A(B[29]), .Y(n147) );
  INVX2 U22 ( .A(B[16]), .Y(n148) );
  INVX2 U23 ( .A(B[15]), .Y(n149) );
  INVX2 U24 ( .A(B[14]), .Y(n150) );
  INVX2 U25 ( .A(B[13]), .Y(n151) );
  INVX2 U26 ( .A(B[12]), .Y(n152) );
  INVX2 U27 ( .A(B[11]), .Y(n153) );
  INVX2 U28 ( .A(B[10]), .Y(n154) );
  INVX2 U29 ( .A(B[9]), .Y(n155) );
  INVX2 U30 ( .A(B[8]), .Y(n156) );
  INVX2 U31 ( .A(B[7]), .Y(n157) );
  INVX2 U32 ( .A(B[6]), .Y(n158) );
  INVX2 U33 ( .A(B[5]), .Y(n159) );
  INVX2 U34 ( .A(B[4]), .Y(n160) );
  INVX2 U35 ( .A(B[3]), .Y(n161) );
  INVX2 U36 ( .A(B[2]), .Y(n162) );
  INVX2 U37 ( .A(B[1]), .Y(n163) );
  INVX2 U38 ( .A(B[0]), .Y(n164) );
  INVX2 U39 ( .A(A[9]), .Y(n165) );
  INVX2 U40 ( .A(A[8]), .Y(n166) );
  INVX2 U41 ( .A(A[30]), .Y(n167) );
  INVX2 U42 ( .A(A[29]), .Y(n168) );
  INVX2 U43 ( .A(A[28]), .Y(n169) );
  INVX2 U44 ( .A(A[27]), .Y(n170) );
  INVX2 U45 ( .A(A[26]), .Y(n171) );
  INVX2 U46 ( .A(A[25]), .Y(n172) );
  INVX2 U47 ( .A(A[24]), .Y(n173) );
  INVX2 U48 ( .A(A[23]), .Y(n174) );
  INVX2 U49 ( .A(A[22]), .Y(n175) );
  INVX2 U50 ( .A(A[21]), .Y(n176) );
  INVX2 U51 ( .A(A[20]), .Y(n177) );
  INVX2 U52 ( .A(A[19]), .Y(n178) );
  INVX2 U53 ( .A(A[18]), .Y(n179) );
  INVX2 U54 ( .A(A[17]), .Y(n180) );
  INVX2 U55 ( .A(A[16]), .Y(n181) );
  INVX2 U56 ( .A(A[15]), .Y(n182) );
  INVX2 U57 ( .A(A[14]), .Y(n183) );
  INVX2 U58 ( .A(A[13]), .Y(n184) );
  INVX2 U59 ( .A(A[12]), .Y(n185) );
  INVX2 U60 ( .A(A[11]), .Y(n186) );
  INVX2 U61 ( .A(A[10]), .Y(n187) );
  INVX2 U62 ( .A(TC), .Y(n188) );
endmodule


module CannyEdge_DW01_add_42 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n141, n142, n143, n144, n145, n146, n147,
         n148, n149;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U31 ( .A(n30), .B(n31), .Y(SUM[9]) );
  NOR2X1 U32 ( .A(n130), .B(n32), .Y(n31) );
  XOR2X1 U33 ( .A(n34), .B(n134), .Y(SUM[8]) );
  NAND2X1 U34 ( .A(n133), .B(n35), .Y(n34) );
  XOR2X1 U35 ( .A(n37), .B(n38), .Y(SUM[7]) );
  XOR2X1 U36 ( .A(n135), .B(B[7]), .Y(n38) );
  OAI21X1 U37 ( .A(B[6]), .B(A[6]), .C(n37), .Y(n39) );
  XOR2X1 U38 ( .A(n40), .B(n41), .Y(SUM[29]) );
  XOR2X1 U39 ( .A(B[29]), .B(A[29]), .Y(n41) );
  OAI21X1 U40 ( .A(n42), .B(n43), .C(n44), .Y(n40) );
  XOR2X1 U41 ( .A(n45), .B(n43), .Y(SUM[28]) );
  AOI21X1 U42 ( .A(n137), .B(n46), .C(n47), .Y(n43) );
  NAND2X1 U43 ( .A(n136), .B(n44), .Y(n45) );
  NAND2X1 U44 ( .A(B[28]), .B(A[28]), .Y(n44) );
  NOR2X1 U45 ( .A(B[28]), .B(A[28]), .Y(n42) );
  XOR2X1 U46 ( .A(n46), .B(n49), .Y(SUM[27]) );
  NOR2X1 U47 ( .A(n47), .B(n48), .Y(n49) );
  NOR2X1 U48 ( .A(B[27]), .B(A[27]), .Y(n48) );
  AND2X1 U49 ( .A(B[27]), .B(A[27]), .Y(n47) );
  OAI21X1 U50 ( .A(n50), .B(n51), .C(n52), .Y(n46) );
  XOR2X1 U51 ( .A(n53), .B(n51), .Y(SUM[26]) );
  AOI21X1 U52 ( .A(n139), .B(n54), .C(n55), .Y(n51) );
  NAND2X1 U53 ( .A(n138), .B(n52), .Y(n53) );
  NAND2X1 U54 ( .A(B[26]), .B(A[26]), .Y(n52) );
  NOR2X1 U55 ( .A(B[26]), .B(A[26]), .Y(n50) );
  XOR2X1 U56 ( .A(n54), .B(n57), .Y(SUM[25]) );
  NOR2X1 U57 ( .A(n55), .B(n56), .Y(n57) );
  NOR2X1 U58 ( .A(B[25]), .B(A[25]), .Y(n56) );
  AND2X1 U59 ( .A(B[25]), .B(A[25]), .Y(n55) );
  OAI21X1 U60 ( .A(n58), .B(n59), .C(n60), .Y(n54) );
  XOR2X1 U61 ( .A(n61), .B(n59), .Y(SUM[24]) );
  AOI21X1 U62 ( .A(n143), .B(n62), .C(n63), .Y(n59) );
  NAND2X1 U63 ( .A(n142), .B(n60), .Y(n61) );
  NAND2X1 U64 ( .A(B[24]), .B(A[24]), .Y(n60) );
  NOR2X1 U65 ( .A(B[24]), .B(A[24]), .Y(n58) );
  XOR2X1 U66 ( .A(n62), .B(n65), .Y(SUM[23]) );
  NOR2X1 U67 ( .A(n63), .B(n64), .Y(n65) );
  NOR2X1 U68 ( .A(B[23]), .B(A[23]), .Y(n64) );
  AND2X1 U69 ( .A(B[23]), .B(A[23]), .Y(n63) );
  OAI21X1 U70 ( .A(n66), .B(n67), .C(n68), .Y(n62) );
  XOR2X1 U71 ( .A(n69), .B(n67), .Y(SUM[22]) );
  AOI21X1 U72 ( .A(n145), .B(n70), .C(n71), .Y(n67) );
  NAND2X1 U73 ( .A(n144), .B(n68), .Y(n69) );
  NAND2X1 U74 ( .A(B[22]), .B(A[22]), .Y(n68) );
  NOR2X1 U75 ( .A(B[22]), .B(A[22]), .Y(n66) );
  XOR2X1 U76 ( .A(n70), .B(n73), .Y(SUM[21]) );
  NOR2X1 U77 ( .A(n71), .B(n72), .Y(n73) );
  NOR2X1 U78 ( .A(B[21]), .B(A[21]), .Y(n72) );
  AND2X1 U79 ( .A(B[21]), .B(A[21]), .Y(n71) );
  OAI21X1 U80 ( .A(n74), .B(n75), .C(n76), .Y(n70) );
  XOR2X1 U81 ( .A(n77), .B(n75), .Y(SUM[20]) );
  AOI21X1 U82 ( .A(n147), .B(n78), .C(n79), .Y(n75) );
  NAND2X1 U83 ( .A(n146), .B(n76), .Y(n77) );
  NAND2X1 U84 ( .A(B[20]), .B(A[20]), .Y(n76) );
  NOR2X1 U85 ( .A(B[20]), .B(A[20]), .Y(n74) );
  XOR2X1 U86 ( .A(n78), .B(n81), .Y(SUM[19]) );
  NOR2X1 U87 ( .A(n79), .B(n80), .Y(n81) );
  NOR2X1 U88 ( .A(B[19]), .B(A[19]), .Y(n80) );
  AND2X1 U89 ( .A(B[19]), .B(A[19]), .Y(n79) );
  OAI21X1 U90 ( .A(n82), .B(n83), .C(n84), .Y(n78) );
  XOR2X1 U91 ( .A(n85), .B(n83), .Y(SUM[18]) );
  AOI21X1 U92 ( .A(n149), .B(n86), .C(n87), .Y(n83) );
  NAND2X1 U93 ( .A(n148), .B(n84), .Y(n85) );
  NAND2X1 U94 ( .A(B[18]), .B(A[18]), .Y(n84) );
  NOR2X1 U95 ( .A(B[18]), .B(A[18]), .Y(n82) );
  XOR2X1 U96 ( .A(n86), .B(n89), .Y(SUM[17]) );
  NOR2X1 U97 ( .A(n87), .B(n88), .Y(n89) );
  NOR2X1 U98 ( .A(B[17]), .B(A[17]), .Y(n88) );
  AND2X1 U99 ( .A(B[17]), .B(A[17]), .Y(n87) );
  OAI21X1 U100 ( .A(n90), .B(n91), .C(n92), .Y(n86) );
  XOR2X1 U101 ( .A(n93), .B(n91), .Y(SUM[16]) );
  AOI21X1 U102 ( .A(n122), .B(n94), .C(n95), .Y(n91) );
  NAND2X1 U103 ( .A(n121), .B(n92), .Y(n93) );
  NAND2X1 U104 ( .A(B[16]), .B(A[16]), .Y(n92) );
  NOR2X1 U105 ( .A(B[16]), .B(A[16]), .Y(n90) );
  XOR2X1 U106 ( .A(n94), .B(n97), .Y(SUM[15]) );
  NOR2X1 U107 ( .A(n95), .B(n96), .Y(n97) );
  NOR2X1 U108 ( .A(B[15]), .B(A[15]), .Y(n96) );
  AND2X1 U109 ( .A(B[15]), .B(A[15]), .Y(n95) );
  OAI21X1 U110 ( .A(n98), .B(n99), .C(n100), .Y(n94) );
  XOR2X1 U111 ( .A(n101), .B(n99), .Y(SUM[14]) );
  AOI21X1 U112 ( .A(n124), .B(n102), .C(n103), .Y(n99) );
  NAND2X1 U113 ( .A(n123), .B(n100), .Y(n101) );
  NAND2X1 U114 ( .A(B[14]), .B(A[14]), .Y(n100) );
  NOR2X1 U115 ( .A(B[14]), .B(A[14]), .Y(n98) );
  XOR2X1 U116 ( .A(n102), .B(n105), .Y(SUM[13]) );
  NOR2X1 U117 ( .A(n103), .B(n104), .Y(n105) );
  NOR2X1 U118 ( .A(B[13]), .B(A[13]), .Y(n104) );
  AND2X1 U119 ( .A(B[13]), .B(A[13]), .Y(n103) );
  OAI21X1 U120 ( .A(n106), .B(n126), .C(n107), .Y(n102) );
  XOR2X1 U121 ( .A(n108), .B(n126), .Y(SUM[12]) );
  OAI21X1 U122 ( .A(n110), .B(n111), .C(n112), .Y(n109) );
  AOI21X1 U123 ( .A(n113), .B(n129), .C(n128), .Y(n111) );
  NAND2X1 U124 ( .A(n125), .B(n107), .Y(n108) );
  NAND2X1 U125 ( .A(B[12]), .B(A[12]), .Y(n107) );
  NOR2X1 U126 ( .A(B[12]), .B(A[12]), .Y(n106) );
  XOR2X1 U127 ( .A(n115), .B(n116), .Y(SUM[11]) );
  NOR2X1 U128 ( .A(n127), .B(n110), .Y(n116) );
  NOR2X1 U129 ( .A(B[11]), .B(A[11]), .Y(n110) );
  NAND2X1 U130 ( .A(B[11]), .B(A[11]), .Y(n112) );
  OAI21X1 U131 ( .A(n117), .B(n131), .C(n114), .Y(n115) );
  XOR2X1 U132 ( .A(n118), .B(n131), .Y(SUM[10]) );
  OAI21X1 U133 ( .A(n132), .B(n32), .C(n33), .Y(n113) );
  NAND2X1 U134 ( .A(B[9]), .B(A[9]), .Y(n33) );
  NOR2X1 U135 ( .A(B[9]), .B(A[9]), .Y(n32) );
  OAI21X1 U136 ( .A(n36), .B(n134), .C(n35), .Y(n30) );
  NAND2X1 U137 ( .A(B[8]), .B(A[8]), .Y(n35) );
  OAI21X1 U138 ( .A(n37), .B(n135), .C(n120), .Y(n119) );
  OAI21X1 U139 ( .A(n141), .B(A[7]), .C(B[7]), .Y(n120) );
  NAND2X1 U140 ( .A(B[6]), .B(A[6]), .Y(n37) );
  NOR2X1 U141 ( .A(B[8]), .B(A[8]), .Y(n36) );
  NAND2X1 U142 ( .A(n129), .B(n114), .Y(n118) );
  NAND2X1 U143 ( .A(B[10]), .B(A[10]), .Y(n114) );
  NOR2X1 U144 ( .A(B[10]), .B(A[10]), .Y(n117) );
  INVX2 U2 ( .A(n90), .Y(n121) );
  INVX2 U3 ( .A(n96), .Y(n122) );
  INVX2 U4 ( .A(n98), .Y(n123) );
  INVX2 U5 ( .A(n104), .Y(n124) );
  INVX2 U6 ( .A(n106), .Y(n125) );
  INVX2 U7 ( .A(n109), .Y(n126) );
  INVX2 U8 ( .A(n112), .Y(n127) );
  INVX2 U9 ( .A(n114), .Y(n128) );
  INVX2 U10 ( .A(n117), .Y(n129) );
  INVX2 U11 ( .A(n33), .Y(n130) );
  INVX2 U12 ( .A(n113), .Y(n131) );
  INVX2 U13 ( .A(n30), .Y(n132) );
  INVX2 U14 ( .A(n36), .Y(n133) );
  INVX2 U15 ( .A(n119), .Y(n134) );
  INVX2 U16 ( .A(A[7]), .Y(n135) );
  INVX2 U17 ( .A(n42), .Y(n136) );
  INVX2 U18 ( .A(n48), .Y(n137) );
  INVX2 U19 ( .A(n50), .Y(n138) );
  INVX2 U20 ( .A(n56), .Y(n139) );
  INVX2 U21 ( .A(n39), .Y(SUM[6]) );
  INVX2 U22 ( .A(n37), .Y(n141) );
  INVX2 U23 ( .A(n58), .Y(n142) );
  INVX2 U24 ( .A(n64), .Y(n143) );
  INVX2 U25 ( .A(n66), .Y(n144) );
  INVX2 U26 ( .A(n72), .Y(n145) );
  INVX2 U27 ( .A(n74), .Y(n146) );
  INVX2 U28 ( .A(n80), .Y(n147) );
  INVX2 U29 ( .A(n82), .Y(n148) );
  INVX2 U30 ( .A(n88), .Y(n149) );
endmodule


module CannyEdge_DW02_mult_20 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][31] , \ab[7][30] , \ab[7][29] , \ab[7][28] , \ab[7][27] ,
         \ab[7][26] , \ab[7][25] , \ab[7][24] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][31] , \ab[6][30] , \ab[6][29] ,
         \ab[6][28] , \ab[6][27] , \ab[6][26] , \ab[6][25] , \ab[6][24] ,
         \ab[6][23] , \ab[6][22] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][31] ,
         \ab[5][30] , \ab[5][29] , \ab[5][28] , \ab[5][27] , \ab[5][26] ,
         \ab[5][25] , \ab[5][24] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][31] , \ab[4][30] , \ab[4][29] , \ab[4][28] ,
         \ab[4][27] , \ab[4][26] , \ab[4][25] , \ab[4][24] , \ab[4][23] ,
         \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][31] , \ab[3][30] ,
         \ab[3][29] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][31] , \ab[2][30] , \ab[2][29] , \ab[2][28] , \ab[2][27] ,
         \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][31] , \ab[1][30] , \ab[1][29] ,
         \ab[1][28] , \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] ,
         \ab[1][23] , \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][31] ,
         \ab[0][30] , \ab[0][29] , \ab[0][28] , \ab[0][27] , \ab[0][26] ,
         \ab[0][25] , \ab[0][24] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[7][31] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][27] , \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][28] , \CARRYB[6][27] ,
         \CARRYB[6][26] , \CARRYB[6][25] , \CARRYB[6][24] , \CARRYB[6][23] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][30] ,
         \CARRYB[5][29] , \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][28] , \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] ,
         \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][30] , \CARRYB[3][29] , \CARRYB[3][28] ,
         \CARRYB[3][27] , \CARRYB[3][26] , \CARRYB[3][25] , \CARRYB[3][24] ,
         \CARRYB[3][23] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][31] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] ,
         \SUMB[6][27] , \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] ,
         \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] ,
         \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] ,
         \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] ,
         \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] ,
         \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] ,
         \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] ,
         \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[30] , n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n111,
         n112, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S14_31_0 ( .A(n120), .B(\CARRYB[7][23] ), .C(\SUMB[7][24] ), .YC(
        \A2[30] ), .YS(\A1[29] ) );
  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S4_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S4_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S4_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S4_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  FAX1 S4_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S4_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S4_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S4_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  FAX1 S4_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S4_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S4_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S4_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  FAX1 S4_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S4_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S4_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S4_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  FAX1 S4_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S4_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S4_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S4_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  FAX1 S4_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S4_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S5_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .C(\ab[6][31] ), .YC(
        \CARRYB[7][30] ), .YS(\SUMB[7][30] ) );
  FAX1 S14_31 ( .A(QA), .B(QB), .C(\ab[7][31] ), .YC(\CARRYB[7][31] ), .YS(
        \SUMB[7][31] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  FAX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  FAX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  FAX1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  FAX1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  FAX1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .C(\ab[5][31] ), .YC(
        \CARRYB[6][30] ), .YS(\SUMB[6][30] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .C(\ab[4][31] ), .YC(
        \CARRYB[5][30] ), .YS(\SUMB[5][30] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .C(\ab[3][31] ), .YC(
        \CARRYB[4][30] ), .YS(\SUMB[4][30] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .C(\ab[2][31] ), .YC(
        \CARRYB[3][30] ), .YS(\SUMB[3][30] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n40), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n39), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n38), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n37), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n36), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n35), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n34), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n33), .C(\SUMB[1][8] ), .YC(\CARRYB[2][7] ), 
        .YS(\SUMB[2][7] ) );
  FAX1 S2_2_8 ( .A(\ab[2][8] ), .B(n32), .C(\SUMB[1][9] ), .YC(\CARRYB[2][8] ), 
        .YS(\SUMB[2][8] ) );
  FAX1 S2_2_9 ( .A(\ab[2][9] ), .B(n31), .C(\SUMB[1][10] ), .YC(\CARRYB[2][9] ), .YS(\SUMB[2][9] ) );
  FAX1 S2_2_10 ( .A(\ab[2][10] ), .B(n30), .C(\SUMB[1][11] ), .YC(
        \CARRYB[2][10] ), .YS(\SUMB[2][10] ) );
  FAX1 S2_2_11 ( .A(\ab[2][11] ), .B(n29), .C(\SUMB[1][12] ), .YC(
        \CARRYB[2][11] ), .YS(\SUMB[2][11] ) );
  FAX1 S2_2_12 ( .A(\ab[2][12] ), .B(n28), .C(\SUMB[1][13] ), .YC(
        \CARRYB[2][12] ), .YS(\SUMB[2][12] ) );
  FAX1 S2_2_13 ( .A(\ab[2][13] ), .B(n27), .C(\SUMB[1][14] ), .YC(
        \CARRYB[2][13] ), .YS(\SUMB[2][13] ) );
  FAX1 S2_2_14 ( .A(\ab[2][14] ), .B(n26), .C(\SUMB[1][15] ), .YC(
        \CARRYB[2][14] ), .YS(\SUMB[2][14] ) );
  FAX1 S2_2_15 ( .A(\ab[2][15] ), .B(n25), .C(\SUMB[1][16] ), .YC(
        \CARRYB[2][15] ), .YS(\SUMB[2][15] ) );
  FAX1 S2_2_16 ( .A(\ab[2][16] ), .B(n24), .C(\SUMB[1][17] ), .YC(
        \CARRYB[2][16] ), .YS(\SUMB[2][16] ) );
  FAX1 S2_2_17 ( .A(\ab[2][17] ), .B(n23), .C(\SUMB[1][18] ), .YC(
        \CARRYB[2][17] ), .YS(\SUMB[2][17] ) );
  FAX1 S2_2_18 ( .A(\ab[2][18] ), .B(n22), .C(\SUMB[1][19] ), .YC(
        \CARRYB[2][18] ), .YS(\SUMB[2][18] ) );
  FAX1 S2_2_19 ( .A(\ab[2][19] ), .B(n21), .C(\SUMB[1][20] ), .YC(
        \CARRYB[2][19] ), .YS(\SUMB[2][19] ) );
  FAX1 S2_2_20 ( .A(\ab[2][20] ), .B(n20), .C(\SUMB[1][21] ), .YC(
        \CARRYB[2][20] ), .YS(\SUMB[2][20] ) );
  FAX1 S2_2_21 ( .A(\ab[2][21] ), .B(n19), .C(\SUMB[1][22] ), .YC(
        \CARRYB[2][21] ), .YS(\SUMB[2][21] ) );
  FAX1 S2_2_22 ( .A(\ab[2][22] ), .B(n18), .C(\SUMB[1][23] ), .YC(
        \CARRYB[2][22] ), .YS(\SUMB[2][22] ) );
  FAX1 S2_2_23 ( .A(\ab[2][23] ), .B(n17), .C(\SUMB[1][24] ), .YC(
        \CARRYB[2][23] ), .YS(\SUMB[2][23] ) );
  FAX1 S2_2_24 ( .A(\ab[2][24] ), .B(n16), .C(\SUMB[1][25] ), .YC(
        \CARRYB[2][24] ), .YS(\SUMB[2][24] ) );
  FAX1 S2_2_25 ( .A(\ab[2][25] ), .B(n15), .C(\SUMB[1][26] ), .YC(
        \CARRYB[2][25] ), .YS(\SUMB[2][25] ) );
  FAX1 S2_2_26 ( .A(\ab[2][26] ), .B(n14), .C(\SUMB[1][27] ), .YC(
        \CARRYB[2][26] ), .YS(\SUMB[2][26] ) );
  FAX1 S2_2_27 ( .A(\ab[2][27] ), .B(n13), .C(\SUMB[1][28] ), .YC(
        \CARRYB[2][27] ), .YS(\SUMB[2][27] ) );
  FAX1 S2_2_28 ( .A(\ab[2][28] ), .B(n12), .C(\SUMB[1][29] ), .YC(
        \CARRYB[2][28] ), .YS(\SUMB[2][28] ) );
  FAX1 S2_2_29 ( .A(\ab[2][29] ), .B(n11), .C(\SUMB[1][30] ), .YC(
        \CARRYB[2][29] ), .YS(\SUMB[2][29] ) );
  FAX1 S3_2_30 ( .A(\ab[2][30] ), .B(n10), .C(\ab[1][31] ), .YC(
        \CARRYB[2][30] ), .YS(\SUMB[2][30] ) );
  AND2X2 U2 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(n3) );
  AND2X2 U3 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(n4) );
  AND2X2 U4 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(n5) );
  AND2X2 U5 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(n6) );
  AND2X2 U6 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(n7) );
  AND2X2 U7 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(n8) );
  AND2X2 U8 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(n9) );
  AND2X2 U9 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Y(n10) );
  AND2X2 U10 ( .A(\ab[0][30] ), .B(\ab[1][29] ), .Y(n11) );
  AND2X2 U11 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Y(n12) );
  AND2X2 U12 ( .A(\ab[0][28] ), .B(\ab[1][27] ), .Y(n13) );
  AND2X2 U13 ( .A(\ab[0][27] ), .B(\ab[1][26] ), .Y(n14) );
  AND2X2 U14 ( .A(\ab[0][26] ), .B(\ab[1][25] ), .Y(n15) );
  AND2X2 U15 ( .A(\ab[0][25] ), .B(\ab[1][24] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[0][24] ), .B(\ab[1][23] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[0][23] ), .B(\ab[1][22] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[0][22] ), .B(\ab[1][21] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Y(n24) );
  AND2X2 U24 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Y(n25) );
  AND2X2 U25 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Y(n26) );
  AND2X2 U26 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Y(n27) );
  AND2X2 U27 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Y(n28) );
  AND2X2 U28 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Y(n29) );
  AND2X2 U29 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Y(n30) );
  AND2X2 U30 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Y(n31) );
  AND2X2 U31 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Y(n36) );
  AND2X2 U36 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Y(n37) );
  AND2X2 U37 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Y(n38) );
  AND2X2 U38 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Y(n39) );
  AND2X2 U39 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n115), .Y(n42) );
  AND2X2 U42 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(n53) );
  AND2X2 U53 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(n54) );
  AND2X2 U54 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(n55) );
  AND2X2 U55 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(n56) );
  AND2X2 U56 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(n57) );
  AND2X2 U57 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(n58) );
  AND2X2 U58 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(n59) );
  AND2X2 U59 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(n60) );
  AND2X2 U60 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(n61) );
  AND2X2 U61 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(n62) );
  AND2X2 U62 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(n63) );
  AND2X2 U63 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(n64) );
  XOR2X1 U67 ( .A(\SUMB[7][0] ), .B(n115), .Y(\A1[5] ) );
  XOR2X1 U68 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  XOR2X1 U69 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  XOR2X1 U70 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  XOR2X1 U71 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  XOR2X1 U72 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  XOR2X1 U73 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  XOR2X1 U74 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  XOR2X1 U75 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  XOR2X1 U76 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  XOR2X1 U77 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  XOR2X1 U78 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  XOR2X1 U79 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  XOR2X1 U80 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  XOR2X1 U81 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  XOR2X1 U82 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  XOR2X1 U83 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  XOR2X1 U84 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  XOR2X1 U85 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  XOR2X1 U86 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  XOR2X1 U87 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  XOR2X1 U88 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  XOR2X1 U89 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  XOR2X1 U90 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  XOR2X1 U91 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  XOR2X1 U92 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  XOR2X1 U93 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  XOR2X1 U94 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  XOR2X1 U95 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  XOR2X1 U96 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  XOR2X1 U97 ( .A(\SUMB[7][31] ), .B(\CARRYB[7][30] ), .Y(\A1[36] ) );
  XOR2X1 U98 ( .A(\CARRYB[7][31] ), .B(TC), .Y(\A1[37] ) );
  XOR2X1 U99 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U100 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U101 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U102 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U103 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U104 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U105 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U106 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Y(\SUMB[1][7] ) );
  XOR2X1 U107 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Y(\SUMB[1][8] ) );
  XOR2X1 U108 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Y(\SUMB[1][9] ) );
  XOR2X1 U109 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Y(\SUMB[1][10] ) );
  XOR2X1 U110 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Y(\SUMB[1][11] ) );
  XOR2X1 U111 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Y(\SUMB[1][12] ) );
  XOR2X1 U112 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Y(\SUMB[1][13] ) );
  XOR2X1 U113 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Y(\SUMB[1][14] ) );
  XOR2X1 U114 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Y(\SUMB[1][15] ) );
  XOR2X1 U115 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Y(\SUMB[1][16] ) );
  XOR2X1 U116 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Y(\SUMB[1][17] ) );
  XOR2X1 U117 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Y(\SUMB[1][18] ) );
  XOR2X1 U118 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Y(\SUMB[1][19] ) );
  XOR2X1 U119 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Y(\SUMB[1][20] ) );
  XOR2X1 U120 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Y(\SUMB[1][21] ) );
  XOR2X1 U121 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Y(\SUMB[1][22] ) );
  XOR2X1 U122 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Y(\SUMB[1][23] ) );
  XOR2X1 U123 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Y(\SUMB[1][24] ) );
  XOR2X1 U124 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Y(\SUMB[1][25] ) );
  XOR2X1 U125 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Y(\SUMB[1][26] ) );
  XOR2X1 U126 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Y(\SUMB[1][27] ) );
  XOR2X1 U127 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Y(\SUMB[1][28] ) );
  XOR2X1 U128 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Y(\SUMB[1][29] ) );
  XOR2X1 U129 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Y(\SUMB[1][30] ) );
  MUX2X1 U170 ( .B(n118), .A(n117), .S(B[9]), .Y(\ab[7][9] ) );
  MUX2X1 U171 ( .B(n118), .A(n117), .S(B[8]), .Y(\ab[7][8] ) );
  MUX2X1 U172 ( .B(n118), .A(n117), .S(B[7]), .Y(\ab[7][7] ) );
  MUX2X1 U173 ( .B(n118), .A(n117), .S(B[6]), .Y(\ab[7][6] ) );
  MUX2X1 U174 ( .B(n118), .A(n117), .S(B[5]), .Y(\ab[7][5] ) );
  MUX2X1 U175 ( .B(n118), .A(n117), .S(B[4]), .Y(\ab[7][4] ) );
  MUX2X1 U176 ( .B(n118), .A(n117), .S(B[3]), .Y(\ab[7][3] ) );
  AND2X1 U177 ( .A(A[7]), .B(B[31]), .Y(\ab[7][31] ) );
  MUX2X1 U178 ( .B(n118), .A(n117), .S(B[30]), .Y(\ab[7][30] ) );
  MUX2X1 U179 ( .B(n118), .A(n117), .S(B[2]), .Y(\ab[7][2] ) );
  MUX2X1 U180 ( .B(n118), .A(n117), .S(B[29]), .Y(\ab[7][29] ) );
  MUX2X1 U181 ( .B(n118), .A(n117), .S(B[28]), .Y(\ab[7][28] ) );
  MUX2X1 U182 ( .B(n118), .A(n117), .S(B[27]), .Y(\ab[7][27] ) );
  MUX2X1 U183 ( .B(n118), .A(n117), .S(B[26]), .Y(\ab[7][26] ) );
  MUX2X1 U184 ( .B(n118), .A(n117), .S(B[25]), .Y(\ab[7][25] ) );
  MUX2X1 U185 ( .B(n118), .A(n117), .S(B[24]), .Y(\ab[7][24] ) );
  MUX2X1 U186 ( .B(n118), .A(n117), .S(B[23]), .Y(\ab[7][23] ) );
  MUX2X1 U187 ( .B(n118), .A(n117), .S(B[22]), .Y(\ab[7][22] ) );
  MUX2X1 U188 ( .B(n118), .A(n117), .S(B[21]), .Y(\ab[7][21] ) );
  MUX2X1 U189 ( .B(n118), .A(n117), .S(B[20]), .Y(\ab[7][20] ) );
  MUX2X1 U190 ( .B(n118), .A(n117), .S(B[1]), .Y(\ab[7][1] ) );
  MUX2X1 U191 ( .B(n118), .A(n117), .S(B[19]), .Y(\ab[7][19] ) );
  MUX2X1 U192 ( .B(n118), .A(n117), .S(B[18]), .Y(\ab[7][18] ) );
  MUX2X1 U193 ( .B(n118), .A(n117), .S(B[17]), .Y(\ab[7][17] ) );
  MUX2X1 U194 ( .B(n118), .A(n117), .S(B[16]), .Y(\ab[7][16] ) );
  MUX2X1 U195 ( .B(n118), .A(n117), .S(B[15]), .Y(\ab[7][15] ) );
  MUX2X1 U196 ( .B(n118), .A(n117), .S(B[14]), .Y(\ab[7][14] ) );
  MUX2X1 U197 ( .B(n118), .A(n117), .S(B[13]), .Y(\ab[7][13] ) );
  MUX2X1 U198 ( .B(n118), .A(n117), .S(B[12]), .Y(\ab[7][12] ) );
  MUX2X1 U199 ( .B(n118), .A(n117), .S(B[11]), .Y(\ab[7][11] ) );
  MUX2X1 U200 ( .B(n118), .A(n117), .S(B[10]), .Y(\ab[7][10] ) );
  MUX2X1 U201 ( .B(n118), .A(n117), .S(B[0]), .Y(\ab[7][0] ) );
  NOR2X1 U203 ( .A(n142), .B(n158), .Y(\ab[6][9] ) );
  NOR2X1 U204 ( .A(n153), .B(n158), .Y(\ab[6][8] ) );
  NOR2X1 U205 ( .A(n152), .B(n158), .Y(\ab[6][7] ) );
  NOR2X1 U206 ( .A(n151), .B(n158), .Y(\ab[6][6] ) );
  NOR2X1 U207 ( .A(n150), .B(n158), .Y(\ab[6][5] ) );
  NOR2X1 U208 ( .A(n149), .B(n158), .Y(\ab[6][4] ) );
  NOR2X1 U209 ( .A(n148), .B(n158), .Y(\ab[6][3] ) );
  MUX2X1 U210 ( .B(n111), .A(n112), .S(A[6]), .Y(\ab[6][31] ) );
  NOR2X1 U211 ( .A(n141), .B(n158), .Y(\ab[6][30] ) );
  NOR2X1 U212 ( .A(n147), .B(n158), .Y(\ab[6][2] ) );
  NOR2X1 U213 ( .A(n140), .B(n158), .Y(\ab[6][29] ) );
  NOR2X1 U214 ( .A(n139), .B(n158), .Y(\ab[6][28] ) );
  NOR2X1 U215 ( .A(n138), .B(n158), .Y(\ab[6][27] ) );
  NOR2X1 U216 ( .A(n137), .B(n158), .Y(\ab[6][26] ) );
  NOR2X1 U217 ( .A(n136), .B(n158), .Y(\ab[6][25] ) );
  NOR2X1 U218 ( .A(n135), .B(n158), .Y(\ab[6][24] ) );
  NOR2X1 U219 ( .A(n134), .B(n158), .Y(\ab[6][23] ) );
  NOR2X1 U220 ( .A(n133), .B(n158), .Y(\ab[6][22] ) );
  NOR2X1 U221 ( .A(n132), .B(n158), .Y(\ab[6][21] ) );
  NOR2X1 U222 ( .A(n131), .B(n158), .Y(\ab[6][20] ) );
  NOR2X1 U223 ( .A(n146), .B(n158), .Y(\ab[6][1] ) );
  NOR2X1 U224 ( .A(n130), .B(n158), .Y(\ab[6][19] ) );
  NOR2X1 U225 ( .A(n129), .B(n158), .Y(\ab[6][18] ) );
  NOR2X1 U226 ( .A(n128), .B(n158), .Y(\ab[6][17] ) );
  NOR2X1 U227 ( .A(n127), .B(n158), .Y(\ab[6][16] ) );
  NOR2X1 U228 ( .A(n126), .B(n158), .Y(\ab[6][15] ) );
  NOR2X1 U229 ( .A(n125), .B(n158), .Y(\ab[6][14] ) );
  NOR2X1 U230 ( .A(n124), .B(n158), .Y(\ab[6][13] ) );
  NOR2X1 U231 ( .A(n123), .B(n158), .Y(\ab[6][12] ) );
  NOR2X1 U232 ( .A(n122), .B(n158), .Y(\ab[6][11] ) );
  NOR2X1 U233 ( .A(n143), .B(n158), .Y(\ab[6][10] ) );
  NOR2X1 U234 ( .A(n145), .B(n158), .Y(\ab[6][0] ) );
  NOR2X1 U235 ( .A(n142), .B(n157), .Y(\ab[5][9] ) );
  NOR2X1 U236 ( .A(n153), .B(n157), .Y(\ab[5][8] ) );
  NOR2X1 U237 ( .A(n152), .B(n157), .Y(\ab[5][7] ) );
  NOR2X1 U238 ( .A(n151), .B(n157), .Y(\ab[5][6] ) );
  NOR2X1 U239 ( .A(n150), .B(n157), .Y(\ab[5][5] ) );
  NOR2X1 U240 ( .A(n149), .B(n157), .Y(\ab[5][4] ) );
  NOR2X1 U241 ( .A(n148), .B(n157), .Y(\ab[5][3] ) );
  MUX2X1 U242 ( .B(n111), .A(n112), .S(A[5]), .Y(\ab[5][31] ) );
  NOR2X1 U243 ( .A(n141), .B(n157), .Y(\ab[5][30] ) );
  NOR2X1 U244 ( .A(n147), .B(n157), .Y(\ab[5][2] ) );
  NOR2X1 U245 ( .A(n140), .B(n157), .Y(\ab[5][29] ) );
  NOR2X1 U246 ( .A(n139), .B(n157), .Y(\ab[5][28] ) );
  NOR2X1 U247 ( .A(n138), .B(n157), .Y(\ab[5][27] ) );
  NOR2X1 U248 ( .A(n137), .B(n157), .Y(\ab[5][26] ) );
  NOR2X1 U249 ( .A(n136), .B(n157), .Y(\ab[5][25] ) );
  NOR2X1 U250 ( .A(n135), .B(n157), .Y(\ab[5][24] ) );
  NOR2X1 U251 ( .A(n134), .B(n157), .Y(\ab[5][23] ) );
  NOR2X1 U252 ( .A(n133), .B(n157), .Y(\ab[5][22] ) );
  NOR2X1 U253 ( .A(n132), .B(n157), .Y(\ab[5][21] ) );
  NOR2X1 U254 ( .A(n131), .B(n157), .Y(\ab[5][20] ) );
  NOR2X1 U255 ( .A(n146), .B(n157), .Y(\ab[5][1] ) );
  NOR2X1 U256 ( .A(n130), .B(n157), .Y(\ab[5][19] ) );
  NOR2X1 U257 ( .A(n129), .B(n157), .Y(\ab[5][18] ) );
  NOR2X1 U258 ( .A(n128), .B(n157), .Y(\ab[5][17] ) );
  NOR2X1 U259 ( .A(n127), .B(n157), .Y(\ab[5][16] ) );
  NOR2X1 U260 ( .A(n126), .B(n157), .Y(\ab[5][15] ) );
  NOR2X1 U261 ( .A(n125), .B(n157), .Y(\ab[5][14] ) );
  NOR2X1 U262 ( .A(n124), .B(n157), .Y(\ab[5][13] ) );
  NOR2X1 U263 ( .A(n123), .B(n157), .Y(\ab[5][12] ) );
  NOR2X1 U264 ( .A(n122), .B(n157), .Y(\ab[5][11] ) );
  NOR2X1 U265 ( .A(n143), .B(n157), .Y(\ab[5][10] ) );
  NOR2X1 U266 ( .A(n145), .B(n157), .Y(\ab[5][0] ) );
  NOR2X1 U267 ( .A(n142), .B(n156), .Y(\ab[4][9] ) );
  NOR2X1 U268 ( .A(n153), .B(n156), .Y(\ab[4][8] ) );
  NOR2X1 U269 ( .A(n152), .B(n156), .Y(\ab[4][7] ) );
  NOR2X1 U270 ( .A(n151), .B(n156), .Y(\ab[4][6] ) );
  NOR2X1 U271 ( .A(n150), .B(n156), .Y(\ab[4][5] ) );
  NOR2X1 U272 ( .A(n149), .B(n156), .Y(\ab[4][4] ) );
  NOR2X1 U273 ( .A(n148), .B(n156), .Y(\ab[4][3] ) );
  MUX2X1 U274 ( .B(n111), .A(n112), .S(A[4]), .Y(\ab[4][31] ) );
  NOR2X1 U275 ( .A(n141), .B(n156), .Y(\ab[4][30] ) );
  NOR2X1 U276 ( .A(n147), .B(n156), .Y(\ab[4][2] ) );
  NOR2X1 U277 ( .A(n140), .B(n156), .Y(\ab[4][29] ) );
  NOR2X1 U278 ( .A(n139), .B(n156), .Y(\ab[4][28] ) );
  NOR2X1 U279 ( .A(n138), .B(n156), .Y(\ab[4][27] ) );
  NOR2X1 U280 ( .A(n137), .B(n156), .Y(\ab[4][26] ) );
  NOR2X1 U281 ( .A(n136), .B(n156), .Y(\ab[4][25] ) );
  NOR2X1 U282 ( .A(n135), .B(n156), .Y(\ab[4][24] ) );
  NOR2X1 U283 ( .A(n134), .B(n156), .Y(\ab[4][23] ) );
  NOR2X1 U284 ( .A(n133), .B(n156), .Y(\ab[4][22] ) );
  NOR2X1 U285 ( .A(n132), .B(n156), .Y(\ab[4][21] ) );
  NOR2X1 U286 ( .A(n131), .B(n156), .Y(\ab[4][20] ) );
  NOR2X1 U287 ( .A(n146), .B(n156), .Y(\ab[4][1] ) );
  NOR2X1 U288 ( .A(n130), .B(n156), .Y(\ab[4][19] ) );
  NOR2X1 U289 ( .A(n129), .B(n156), .Y(\ab[4][18] ) );
  NOR2X1 U290 ( .A(n128), .B(n156), .Y(\ab[4][17] ) );
  NOR2X1 U291 ( .A(n127), .B(n156), .Y(\ab[4][16] ) );
  NOR2X1 U292 ( .A(n126), .B(n156), .Y(\ab[4][15] ) );
  NOR2X1 U293 ( .A(n125), .B(n156), .Y(\ab[4][14] ) );
  NOR2X1 U294 ( .A(n124), .B(n156), .Y(\ab[4][13] ) );
  NOR2X1 U295 ( .A(n123), .B(n156), .Y(\ab[4][12] ) );
  NOR2X1 U296 ( .A(n122), .B(n156), .Y(\ab[4][11] ) );
  NOR2X1 U297 ( .A(n143), .B(n156), .Y(\ab[4][10] ) );
  NOR2X1 U298 ( .A(n145), .B(n156), .Y(\ab[4][0] ) );
  NOR2X1 U299 ( .A(n142), .B(n155), .Y(\ab[3][9] ) );
  NOR2X1 U300 ( .A(n153), .B(n155), .Y(\ab[3][8] ) );
  NOR2X1 U301 ( .A(n152), .B(n155), .Y(\ab[3][7] ) );
  NOR2X1 U302 ( .A(n151), .B(n155), .Y(\ab[3][6] ) );
  NOR2X1 U303 ( .A(n150), .B(n155), .Y(\ab[3][5] ) );
  NOR2X1 U304 ( .A(n149), .B(n155), .Y(\ab[3][4] ) );
  NOR2X1 U305 ( .A(n148), .B(n155), .Y(\ab[3][3] ) );
  MUX2X1 U306 ( .B(n111), .A(n112), .S(A[3]), .Y(\ab[3][31] ) );
  NOR2X1 U307 ( .A(n141), .B(n155), .Y(\ab[3][30] ) );
  NOR2X1 U308 ( .A(n147), .B(n155), .Y(\ab[3][2] ) );
  NOR2X1 U309 ( .A(n140), .B(n155), .Y(\ab[3][29] ) );
  NOR2X1 U310 ( .A(n139), .B(n155), .Y(\ab[3][28] ) );
  NOR2X1 U311 ( .A(n138), .B(n155), .Y(\ab[3][27] ) );
  NOR2X1 U312 ( .A(n137), .B(n155), .Y(\ab[3][26] ) );
  NOR2X1 U313 ( .A(n136), .B(n155), .Y(\ab[3][25] ) );
  NOR2X1 U314 ( .A(n135), .B(n155), .Y(\ab[3][24] ) );
  NOR2X1 U315 ( .A(n134), .B(n155), .Y(\ab[3][23] ) );
  NOR2X1 U316 ( .A(n133), .B(n155), .Y(\ab[3][22] ) );
  NOR2X1 U317 ( .A(n132), .B(n155), .Y(\ab[3][21] ) );
  NOR2X1 U318 ( .A(n131), .B(n155), .Y(\ab[3][20] ) );
  NOR2X1 U319 ( .A(n146), .B(n155), .Y(\ab[3][1] ) );
  NOR2X1 U320 ( .A(n130), .B(n155), .Y(\ab[3][19] ) );
  NOR2X1 U321 ( .A(n129), .B(n155), .Y(\ab[3][18] ) );
  NOR2X1 U322 ( .A(n128), .B(n155), .Y(\ab[3][17] ) );
  NOR2X1 U323 ( .A(n127), .B(n155), .Y(\ab[3][16] ) );
  NOR2X1 U324 ( .A(n126), .B(n155), .Y(\ab[3][15] ) );
  NOR2X1 U325 ( .A(n125), .B(n155), .Y(\ab[3][14] ) );
  NOR2X1 U326 ( .A(n124), .B(n155), .Y(\ab[3][13] ) );
  NOR2X1 U327 ( .A(n123), .B(n155), .Y(\ab[3][12] ) );
  NOR2X1 U328 ( .A(n122), .B(n155), .Y(\ab[3][11] ) );
  NOR2X1 U329 ( .A(n143), .B(n155), .Y(\ab[3][10] ) );
  NOR2X1 U330 ( .A(n145), .B(n155), .Y(\ab[3][0] ) );
  NOR2X1 U331 ( .A(n142), .B(n144), .Y(\ab[2][9] ) );
  NOR2X1 U332 ( .A(n153), .B(n144), .Y(\ab[2][8] ) );
  NOR2X1 U333 ( .A(n152), .B(n144), .Y(\ab[2][7] ) );
  NOR2X1 U334 ( .A(n151), .B(n144), .Y(\ab[2][6] ) );
  NOR2X1 U335 ( .A(n150), .B(n144), .Y(\ab[2][5] ) );
  NOR2X1 U336 ( .A(n149), .B(n144), .Y(\ab[2][4] ) );
  NOR2X1 U337 ( .A(n148), .B(n144), .Y(\ab[2][3] ) );
  MUX2X1 U338 ( .B(n111), .A(n112), .S(A[2]), .Y(\ab[2][31] ) );
  NOR2X1 U339 ( .A(n141), .B(n144), .Y(\ab[2][30] ) );
  NOR2X1 U340 ( .A(n147), .B(n144), .Y(\ab[2][2] ) );
  NOR2X1 U341 ( .A(n140), .B(n144), .Y(\ab[2][29] ) );
  NOR2X1 U342 ( .A(n139), .B(n144), .Y(\ab[2][28] ) );
  NOR2X1 U343 ( .A(n138), .B(n144), .Y(\ab[2][27] ) );
  NOR2X1 U344 ( .A(n137), .B(n144), .Y(\ab[2][26] ) );
  NOR2X1 U345 ( .A(n136), .B(n144), .Y(\ab[2][25] ) );
  NOR2X1 U346 ( .A(n135), .B(n144), .Y(\ab[2][24] ) );
  NOR2X1 U347 ( .A(n134), .B(n144), .Y(\ab[2][23] ) );
  NOR2X1 U348 ( .A(n133), .B(n144), .Y(\ab[2][22] ) );
  NOR2X1 U349 ( .A(n132), .B(n144), .Y(\ab[2][21] ) );
  NOR2X1 U350 ( .A(n131), .B(n144), .Y(\ab[2][20] ) );
  NOR2X1 U351 ( .A(n146), .B(n144), .Y(\ab[2][1] ) );
  NOR2X1 U352 ( .A(n130), .B(n144), .Y(\ab[2][19] ) );
  NOR2X1 U353 ( .A(n129), .B(n144), .Y(\ab[2][18] ) );
  NOR2X1 U354 ( .A(n128), .B(n144), .Y(\ab[2][17] ) );
  NOR2X1 U355 ( .A(n127), .B(n144), .Y(\ab[2][16] ) );
  NOR2X1 U356 ( .A(n126), .B(n144), .Y(\ab[2][15] ) );
  NOR2X1 U357 ( .A(n125), .B(n144), .Y(\ab[2][14] ) );
  NOR2X1 U358 ( .A(n124), .B(n144), .Y(\ab[2][13] ) );
  NOR2X1 U359 ( .A(n123), .B(n144), .Y(\ab[2][12] ) );
  NOR2X1 U360 ( .A(n122), .B(n144), .Y(\ab[2][11] ) );
  NOR2X1 U361 ( .A(n143), .B(n144), .Y(\ab[2][10] ) );
  NOR2X1 U362 ( .A(n145), .B(n144), .Y(\ab[2][0] ) );
  NOR2X1 U363 ( .A(n142), .B(n154), .Y(\ab[1][9] ) );
  NOR2X1 U364 ( .A(n153), .B(n154), .Y(\ab[1][8] ) );
  NOR2X1 U365 ( .A(n152), .B(n154), .Y(\ab[1][7] ) );
  NOR2X1 U366 ( .A(n151), .B(n154), .Y(\ab[1][6] ) );
  NOR2X1 U367 ( .A(n150), .B(n154), .Y(\ab[1][5] ) );
  NOR2X1 U368 ( .A(n149), .B(n154), .Y(\ab[1][4] ) );
  NOR2X1 U369 ( .A(n148), .B(n154), .Y(\ab[1][3] ) );
  MUX2X1 U370 ( .B(n111), .A(n112), .S(A[1]), .Y(\ab[1][31] ) );
  NOR2X1 U371 ( .A(n141), .B(n154), .Y(\ab[1][30] ) );
  NOR2X1 U372 ( .A(n147), .B(n154), .Y(\ab[1][2] ) );
  NOR2X1 U373 ( .A(n140), .B(n154), .Y(\ab[1][29] ) );
  NOR2X1 U374 ( .A(n139), .B(n154), .Y(\ab[1][28] ) );
  NOR2X1 U375 ( .A(n138), .B(n154), .Y(\ab[1][27] ) );
  NOR2X1 U376 ( .A(n137), .B(n154), .Y(\ab[1][26] ) );
  NOR2X1 U377 ( .A(n136), .B(n154), .Y(\ab[1][25] ) );
  NOR2X1 U378 ( .A(n135), .B(n154), .Y(\ab[1][24] ) );
  NOR2X1 U379 ( .A(n134), .B(n154), .Y(\ab[1][23] ) );
  NOR2X1 U380 ( .A(n133), .B(n154), .Y(\ab[1][22] ) );
  NOR2X1 U381 ( .A(n132), .B(n154), .Y(\ab[1][21] ) );
  NOR2X1 U382 ( .A(n131), .B(n154), .Y(\ab[1][20] ) );
  NOR2X1 U383 ( .A(n146), .B(n154), .Y(\ab[1][1] ) );
  NOR2X1 U384 ( .A(n130), .B(n154), .Y(\ab[1][19] ) );
  NOR2X1 U385 ( .A(n129), .B(n154), .Y(\ab[1][18] ) );
  NOR2X1 U386 ( .A(n128), .B(n154), .Y(\ab[1][17] ) );
  NOR2X1 U387 ( .A(n127), .B(n154), .Y(\ab[1][16] ) );
  NOR2X1 U388 ( .A(n126), .B(n154), .Y(\ab[1][15] ) );
  NOR2X1 U389 ( .A(n125), .B(n154), .Y(\ab[1][14] ) );
  NOR2X1 U390 ( .A(n124), .B(n154), .Y(\ab[1][13] ) );
  NOR2X1 U391 ( .A(n123), .B(n154), .Y(\ab[1][12] ) );
  NOR2X1 U392 ( .A(n122), .B(n154), .Y(\ab[1][11] ) );
  NOR2X1 U393 ( .A(n143), .B(n154), .Y(\ab[1][10] ) );
  NOR2X1 U394 ( .A(n145), .B(n154), .Y(\ab[1][0] ) );
  NOR2X1 U395 ( .A(n142), .B(n121), .Y(\ab[0][9] ) );
  NOR2X1 U396 ( .A(n153), .B(n121), .Y(\ab[0][8] ) );
  NOR2X1 U397 ( .A(n152), .B(n121), .Y(\ab[0][7] ) );
  NOR2X1 U398 ( .A(n151), .B(n121), .Y(\ab[0][6] ) );
  NOR2X1 U399 ( .A(n150), .B(n121), .Y(\ab[0][5] ) );
  NOR2X1 U400 ( .A(n149), .B(n121), .Y(\ab[0][4] ) );
  NOR2X1 U401 ( .A(n148), .B(n121), .Y(\ab[0][3] ) );
  MUX2X1 U402 ( .B(n111), .A(n112), .S(A[0]), .Y(\ab[0][31] ) );
  NAND2X1 U403 ( .A(B[31]), .B(n119), .Y(n112) );
  NOR2X1 U404 ( .A(n141), .B(n121), .Y(\ab[0][30] ) );
  NOR2X1 U405 ( .A(n147), .B(n121), .Y(\ab[0][2] ) );
  NOR2X1 U406 ( .A(n140), .B(n121), .Y(\ab[0][29] ) );
  NOR2X1 U407 ( .A(n139), .B(n121), .Y(\ab[0][28] ) );
  NOR2X1 U408 ( .A(n138), .B(n121), .Y(\ab[0][27] ) );
  NOR2X1 U409 ( .A(n137), .B(n121), .Y(\ab[0][26] ) );
  NOR2X1 U410 ( .A(n136), .B(n121), .Y(\ab[0][25] ) );
  NOR2X1 U411 ( .A(n135), .B(n121), .Y(\ab[0][24] ) );
  NOR2X1 U412 ( .A(n134), .B(n121), .Y(\ab[0][23] ) );
  NOR2X1 U413 ( .A(n133), .B(n121), .Y(\ab[0][22] ) );
  NOR2X1 U414 ( .A(n132), .B(n121), .Y(\ab[0][21] ) );
  NOR2X1 U415 ( .A(n131), .B(n121), .Y(\ab[0][20] ) );
  NOR2X1 U416 ( .A(n146), .B(n121), .Y(\ab[0][1] ) );
  NOR2X1 U417 ( .A(n130), .B(n121), .Y(\ab[0][19] ) );
  NOR2X1 U418 ( .A(n129), .B(n121), .Y(\ab[0][18] ) );
  NOR2X1 U419 ( .A(n128), .B(n121), .Y(\ab[0][17] ) );
  NOR2X1 U420 ( .A(n127), .B(n121), .Y(\ab[0][16] ) );
  NOR2X1 U421 ( .A(n126), .B(n121), .Y(\ab[0][15] ) );
  NOR2X1 U422 ( .A(n125), .B(n121), .Y(\ab[0][14] ) );
  NOR2X1 U423 ( .A(n124), .B(n121), .Y(\ab[0][13] ) );
  NOR2X1 U424 ( .A(n123), .B(n121), .Y(\ab[0][12] ) );
  NOR2X1 U425 ( .A(n122), .B(n121), .Y(\ab[0][11] ) );
  NOR2X1 U426 ( .A(n143), .B(n121), .Y(\ab[0][10] ) );
  NAND2X1 U427 ( .A(B[31]), .B(TC), .Y(n111) );
  NOR2X1 U429 ( .A(B[31]), .B(n119), .Y(QB) );
  NOR2X1 U430 ( .A(A[7]), .B(n119), .Y(QA) );
  NOR2X1 U431 ( .A(n145), .B(n121), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_42 FS_1 ( .A({\A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n9, n8, n7, 
        n6, n5, n4, n3, \A2[30] , n43, n52, n44, n53, n45, n54, n46, n55, n47, 
        n56, n48, n57, n49, n63, n51, n64, n50, n58, n59, n62, n60, n61, n41, 
        n42, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  AND2X2 U66 ( .A(TC), .B(A[7]), .Y(n115) );
  AND2X2 U130 ( .A(A[7]), .B(n119), .Y(n116) );
  INVX2 U131 ( .A(n116), .Y(n117) );
  INVX2 U132 ( .A(n115), .Y(n118) );
  INVX2 U133 ( .A(TC), .Y(n119) );
  INVX2 U134 ( .A(n111), .Y(n120) );
  INVX2 U135 ( .A(A[0]), .Y(n121) );
  INVX2 U136 ( .A(B[11]), .Y(n122) );
  INVX2 U137 ( .A(B[12]), .Y(n123) );
  INVX2 U138 ( .A(B[13]), .Y(n124) );
  INVX2 U139 ( .A(B[14]), .Y(n125) );
  INVX2 U140 ( .A(B[15]), .Y(n126) );
  INVX2 U141 ( .A(B[16]), .Y(n127) );
  INVX2 U142 ( .A(B[17]), .Y(n128) );
  INVX2 U143 ( .A(B[18]), .Y(n129) );
  INVX2 U144 ( .A(B[19]), .Y(n130) );
  INVX2 U145 ( .A(B[20]), .Y(n131) );
  INVX2 U146 ( .A(B[21]), .Y(n132) );
  INVX2 U147 ( .A(B[22]), .Y(n133) );
  INVX2 U148 ( .A(B[23]), .Y(n134) );
  INVX2 U149 ( .A(B[24]), .Y(n135) );
  INVX2 U150 ( .A(B[25]), .Y(n136) );
  INVX2 U151 ( .A(B[26]), .Y(n137) );
  INVX2 U152 ( .A(B[27]), .Y(n138) );
  INVX2 U153 ( .A(B[28]), .Y(n139) );
  INVX2 U154 ( .A(B[29]), .Y(n140) );
  INVX2 U155 ( .A(B[30]), .Y(n141) );
  INVX2 U156 ( .A(B[9]), .Y(n142) );
  INVX2 U157 ( .A(B[10]), .Y(n143) );
  INVX2 U158 ( .A(A[2]), .Y(n144) );
  INVX2 U159 ( .A(B[0]), .Y(n145) );
  INVX2 U160 ( .A(B[1]), .Y(n146) );
  INVX2 U161 ( .A(B[2]), .Y(n147) );
  INVX2 U162 ( .A(B[3]), .Y(n148) );
  INVX2 U163 ( .A(B[4]), .Y(n149) );
  INVX2 U164 ( .A(B[5]), .Y(n150) );
  INVX2 U165 ( .A(B[6]), .Y(n151) );
  INVX2 U166 ( .A(B[7]), .Y(n152) );
  INVX2 U167 ( .A(B[8]), .Y(n153) );
  INVX2 U168 ( .A(A[1]), .Y(n154) );
  INVX2 U169 ( .A(A[3]), .Y(n155) );
  INVX2 U202 ( .A(A[4]), .Y(n156) );
  INVX2 U428 ( .A(A[5]), .Y(n157) );
  INVX2 U432 ( .A(A[6]), .Y(n158) );
endmodule


module CannyEdge_DW02_mult_21 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] ,
         \SUMB[7][1] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] ,
         \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[9] , \A1[8] , \A1[7] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n60, n61, n62, n63;
  assign \ab[2][7]  = B[7];
  assign \ab[2][6]  = B[6];
  assign \ab[2][5]  = B[5];
  assign \ab[2][4]  = B[4];
  assign \ab[2][3]  = B[3];
  assign \ab[2][2]  = B[2];
  assign \ab[2][1]  = B[1];
  assign PRODUCT[0] = \ab[2][0] ;
  assign \ab[2][0]  = B[0];

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n17), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(PRODUCT[2]) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n20), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n18), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n19), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n16), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n22), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n21), .C(\ab[2][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U2 ( .A(n61), .B(n23), .Y(PRODUCT[9]) );
  AND2X2 U3 ( .A(n28), .B(\SUMB[5][5] ), .Y(n4) );
  AND2X2 U4 ( .A(n29), .B(\SUMB[6][1] ), .Y(n5) );
  AND2X2 U5 ( .A(n32), .B(\SUMB[5][4] ), .Y(n6) );
  AND2X2 U6 ( .A(n33), .B(\SUMB[3][1] ), .Y(n7) );
  AND2X2 U7 ( .A(n34), .B(\SUMB[3][2] ), .Y(n8) );
  AND2X2 U8 ( .A(n38), .B(\SUMB[3][3] ), .Y(n9) );
  AND2X2 U9 ( .A(n35), .B(\SUMB[3][4] ), .Y(n10) );
  AND2X2 U10 ( .A(n36), .B(\SUMB[3][5] ), .Y(n11) );
  AND2X2 U11 ( .A(n37), .B(\SUMB[3][6] ), .Y(n12) );
  AND2X2 U12 ( .A(n30), .B(\SUMB[6][2] ), .Y(n13) );
  AND2X2 U13 ( .A(n31), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(\SUMB[7][4] ), .B(n24), .Y(n15) );
  AND2X2 U15 ( .A(\ab[2][5] ), .B(\ab[2][4] ), .Y(n16) );
  AND2X2 U16 ( .A(\ab[2][1] ), .B(\ab[2][0] ), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][3] ), .B(\ab[2][2] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][4] ), .B(\ab[2][3] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][2] ), .B(\ab[2][1] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][7] ), .B(\ab[2][6] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][6] ), .B(\ab[2][5] ), .Y(n22) );
  AND2X2 U22 ( .A(n5), .B(\SUMB[7][1] ), .Y(n23) );
  AND2X2 U23 ( .A(n6), .B(\SUMB[6][4] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[4][1] ), .Y(n25) );
  AND2X2 U25 ( .A(n8), .B(\SUMB[4][2] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[4][3] ), .Y(n27) );
  AND2X2 U27 ( .A(n11), .B(\SUMB[4][5] ), .Y(n28) );
  AND2X2 U28 ( .A(n25), .B(\SUMB[5][1] ), .Y(n29) );
  AND2X2 U29 ( .A(n26), .B(\SUMB[5][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n27), .B(\SUMB[5][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n10), .B(\SUMB[4][4] ), .Y(n32) );
  AND2X2 U32 ( .A(\CARRYB[2][0] ), .B(\SUMB[2][1] ), .Y(n33) );
  AND2X2 U33 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n34) );
  AND2X2 U34 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n35) );
  AND2X2 U35 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n36) );
  AND2X2 U36 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n37) );
  AND2X2 U37 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n38) );
  AND2X2 U38 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n39) );
  AND2X2 U39 ( .A(n12), .B(n39), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[7][3] ), .B(n14), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][2] ), .B(n13), .Y(n42) );
  AND2X2 U42 ( .A(n4), .B(n40), .Y(n43) );
  XOR2X1 U43 ( .A(\SUMB[7][1] ), .B(n5), .Y(PRODUCT[8]) );
  XOR2X1 U44 ( .A(\SUMB[7][2] ), .B(n13), .Y(\A1[7] ) );
  XOR2X1 U45 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U46 ( .A(\SUMB[7][4] ), .B(n24), .Y(\A1[9] ) );
  XOR2X1 U47 ( .A(\ab[2][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U48 ( .A(\ab[2][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U49 ( .A(\ab[2][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U50 ( .A(\ab[2][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U51 ( .A(\ab[2][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U52 ( .A(\ab[2][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U53 ( .A(\ab[2][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U54 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(PRODUCT[3]) );
  XOR2X1 U55 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U57 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U58 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U59 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U60 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n33), .Y(PRODUCT[4]) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n34), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n38), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n35), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n36), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(\SUMB[3][6] ), .B(n37), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n7), .Y(PRODUCT[5]) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n8), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n9), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n10), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n11), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n39), .B(n12), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n25), .Y(PRODUCT[6]) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n26), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n27), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n32), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n28), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(\SUMB[6][1] ), .B(n29), .Y(PRODUCT[7]) );
  XOR2X1 U79 ( .A(\SUMB[6][2] ), .B(n30), .Y(\SUMB[7][1] ) );
  XOR2X1 U80 ( .A(\SUMB[6][3] ), .B(n31), .Y(\SUMB[7][2] ) );
  XOR2X1 U81 ( .A(\SUMB[6][4] ), .B(n6), .Y(\SUMB[7][3] ) );
  XOR2X1 U82 ( .A(n40), .B(n4), .Y(\SUMB[7][4] ) );
  NOR2X1 U83 ( .A(n15), .B(n43), .Y(n48) );
  NAND2X1 U84 ( .A(n15), .B(n43), .Y(n46) );
  NAND2X1 U85 ( .A(n63), .B(n46), .Y(n45) );
  NOR2X1 U86 ( .A(n42), .B(\A1[8] ), .Y(n49) );
  NAND2X1 U87 ( .A(n42), .B(\A1[8] ), .Y(n50) );
  OAI21X1 U88 ( .A(n44), .B(n49), .C(n50), .Y(n55) );
  NOR2X1 U89 ( .A(n41), .B(\A1[9] ), .Y(n52) );
  AND2X1 U90 ( .A(n41), .B(\A1[9] ), .Y(n53) );
  AOI21X1 U91 ( .A(n55), .B(n62), .C(n53), .Y(n47) );
  XOR2X1 U92 ( .A(n45), .B(n47), .Y(PRODUCT[12]) );
  OAI21X1 U93 ( .A(n48), .B(n47), .C(n46), .Y(PRODUCT[13]) );
  NAND2X1 U94 ( .A(n60), .B(n50), .Y(n51) );
  XOR2X1 U95 ( .A(n51), .B(n44), .Y(PRODUCT[10]) );
  NOR2X1 U96 ( .A(n53), .B(n52), .Y(n54) );
  XOR2X1 U97 ( .A(n55), .B(n54), .Y(PRODUCT[11]) );
  NAND2X1 U98 ( .A(\A1[7] ), .B(n23), .Y(n44) );
  INVX2 U99 ( .A(n49), .Y(n60) );
  INVX2 U100 ( .A(\A1[7] ), .Y(n61) );
  INVX2 U101 ( .A(n52), .Y(n62) );
  INVX2 U102 ( .A(n48), .Y(n63) );
endmodule


module CannyEdge_DW01_cmp2_5 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180;

  MUX2X1 U60 ( .B(n60), .A(n61), .S(B[31]), .Y(LT_LE) );
  MUX2X1 U61 ( .B(n158), .A(n62), .S(A[31]), .Y(n61) );
  NAND2X1 U62 ( .A(A[30]), .B(n63), .Y(n62) );
  MUX2X1 U63 ( .B(n122), .A(TC), .S(A[31]), .Y(n60) );
  OAI21X1 U64 ( .A(B[31]), .B(n178), .C(n64), .Y(n63) );
  AOI21X1 U65 ( .A(A[29]), .B(n137), .C(n65), .Y(n64) );
  AOI21X1 U66 ( .A(B[29]), .B(n177), .C(n66), .Y(n65) );
  OAI21X1 U67 ( .A(A[28]), .B(n138), .C(n67), .Y(n66) );
  OAI21X1 U68 ( .A(B[28]), .B(n176), .C(n68), .Y(n67) );
  AOI21X1 U69 ( .A(A[27]), .B(n139), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(B[27]), .B(n175), .C(n70), .Y(n69) );
  OAI21X1 U71 ( .A(A[26]), .B(n140), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(B[26]), .B(n174), .C(n72), .Y(n71) );
  AOI21X1 U73 ( .A(A[25]), .B(n141), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(B[25]), .B(n173), .C(n74), .Y(n73) );
  OAI21X1 U75 ( .A(A[24]), .B(n142), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(B[24]), .B(n172), .C(n76), .Y(n75) );
  AOI21X1 U77 ( .A(A[23]), .B(n143), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(B[23]), .B(n171), .C(n78), .Y(n77) );
  OAI21X1 U79 ( .A(A[22]), .B(n144), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(B[22]), .B(n170), .C(n80), .Y(n79) );
  AOI21X1 U81 ( .A(A[21]), .B(n145), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(B[21]), .B(n169), .C(n82), .Y(n81) );
  OAI21X1 U83 ( .A(A[20]), .B(n146), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(B[20]), .B(n168), .C(n84), .Y(n83) );
  AOI21X1 U85 ( .A(A[19]), .B(n147), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(B[19]), .B(n167), .C(n86), .Y(n85) );
  OAI21X1 U87 ( .A(A[18]), .B(n148), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(B[18]), .B(n166), .C(n88), .Y(n87) );
  AOI21X1 U89 ( .A(A[17]), .B(n149), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(B[17]), .B(n165), .C(n90), .Y(n89) );
  OAI21X1 U91 ( .A(A[16]), .B(n150), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(B[16]), .B(n164), .C(n92), .Y(n91) );
  AOI21X1 U93 ( .A(A[15]), .B(n151), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(B[15]), .B(n163), .C(n94), .Y(n93) );
  OAI21X1 U95 ( .A(A[14]), .B(n152), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(B[14]), .B(n162), .C(n96), .Y(n95) );
  AOI21X1 U97 ( .A(A[13]), .B(n153), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(B[13]), .B(n161), .C(n98), .Y(n97) );
  OAI21X1 U99 ( .A(A[12]), .B(n154), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(B[12]), .B(n160), .C(n100), .Y(n99) );
  AOI21X1 U101 ( .A(A[11]), .B(n155), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(B[11]), .B(n159), .C(n102), .Y(n101) );
  OAI21X1 U103 ( .A(A[10]), .B(n156), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(B[9]), .B(n180), .C(n104), .Y(n103) );
  AOI21X1 U105 ( .A(A[10]), .B(n156), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(B[9]), .B(n180), .C(n106), .Y(n105) );
  OAI21X1 U107 ( .A(A[8]), .B(n157), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(B[8]), .B(n179), .C(n108), .Y(n107) );
  AOI21X1 U109 ( .A(A[7]), .B(n126), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(B[7]), .B(n136), .C(n110), .Y(n109) );
  OAI21X1 U111 ( .A(A[6]), .B(n125), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(B[6]), .B(n135), .C(n112), .Y(n111) );
  AOI21X1 U113 ( .A(A[5]), .B(n124), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(B[5]), .B(n134), .C(n114), .Y(n113) );
  OAI21X1 U115 ( .A(A[4]), .B(n123), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(B[4]), .B(n133), .C(n116), .Y(n115) );
  AOI21X1 U117 ( .A(A[3]), .B(n129), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(B[3]), .B(n130), .C(n118), .Y(n117) );
  OAI21X1 U119 ( .A(A[2]), .B(n128), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(B[2]), .B(n132), .C(n120), .Y(n119) );
  AOI22X1 U121 ( .A(n121), .B(A[0]), .C(A[1]), .D(n127), .Y(n120) );
  AOI21X1 U122 ( .A(B[1]), .B(n131), .C(B[0]), .Y(n121) );
  INVX2 U1 ( .A(n63), .Y(n122) );
  INVX2 U2 ( .A(B[4]), .Y(n123) );
  INVX2 U3 ( .A(B[5]), .Y(n124) );
  INVX2 U4 ( .A(B[6]), .Y(n125) );
  INVX2 U5 ( .A(B[7]), .Y(n126) );
  INVX2 U6 ( .A(B[1]), .Y(n127) );
  INVX2 U7 ( .A(B[2]), .Y(n128) );
  INVX2 U8 ( .A(B[3]), .Y(n129) );
  INVX2 U9 ( .A(A[3]), .Y(n130) );
  INVX2 U10 ( .A(A[1]), .Y(n131) );
  INVX2 U11 ( .A(A[2]), .Y(n132) );
  INVX2 U12 ( .A(A[4]), .Y(n133) );
  INVX2 U13 ( .A(A[5]), .Y(n134) );
  INVX2 U14 ( .A(A[6]), .Y(n135) );
  INVX2 U15 ( .A(A[7]), .Y(n136) );
  INVX2 U16 ( .A(B[29]), .Y(n137) );
  INVX2 U17 ( .A(B[28]), .Y(n138) );
  INVX2 U18 ( .A(B[27]), .Y(n139) );
  INVX2 U19 ( .A(B[26]), .Y(n140) );
  INVX2 U20 ( .A(B[25]), .Y(n141) );
  INVX2 U21 ( .A(B[24]), .Y(n142) );
  INVX2 U22 ( .A(B[23]), .Y(n143) );
  INVX2 U23 ( .A(B[22]), .Y(n144) );
  INVX2 U24 ( .A(B[21]), .Y(n145) );
  INVX2 U25 ( .A(B[20]), .Y(n146) );
  INVX2 U26 ( .A(B[19]), .Y(n147) );
  INVX2 U27 ( .A(B[18]), .Y(n148) );
  INVX2 U28 ( .A(B[17]), .Y(n149) );
  INVX2 U29 ( .A(B[16]), .Y(n150) );
  INVX2 U30 ( .A(B[15]), .Y(n151) );
  INVX2 U31 ( .A(B[14]), .Y(n152) );
  INVX2 U32 ( .A(B[13]), .Y(n153) );
  INVX2 U33 ( .A(B[12]), .Y(n154) );
  INVX2 U34 ( .A(B[11]), .Y(n155) );
  INVX2 U35 ( .A(B[10]), .Y(n156) );
  INVX2 U36 ( .A(B[8]), .Y(n157) );
  INVX2 U37 ( .A(TC), .Y(n158) );
  INVX2 U38 ( .A(A[11]), .Y(n159) );
  INVX2 U39 ( .A(A[12]), .Y(n160) );
  INVX2 U40 ( .A(A[13]), .Y(n161) );
  INVX2 U41 ( .A(A[14]), .Y(n162) );
  INVX2 U42 ( .A(A[15]), .Y(n163) );
  INVX2 U43 ( .A(A[16]), .Y(n164) );
  INVX2 U44 ( .A(A[17]), .Y(n165) );
  INVX2 U45 ( .A(A[18]), .Y(n166) );
  INVX2 U46 ( .A(A[19]), .Y(n167) );
  INVX2 U47 ( .A(A[20]), .Y(n168) );
  INVX2 U48 ( .A(A[21]), .Y(n169) );
  INVX2 U49 ( .A(A[22]), .Y(n170) );
  INVX2 U50 ( .A(A[23]), .Y(n171) );
  INVX2 U51 ( .A(A[24]), .Y(n172) );
  INVX2 U52 ( .A(A[25]), .Y(n173) );
  INVX2 U53 ( .A(A[26]), .Y(n174) );
  INVX2 U54 ( .A(A[27]), .Y(n175) );
  INVX2 U55 ( .A(A[28]), .Y(n176) );
  INVX2 U56 ( .A(A[29]), .Y(n177) );
  INVX2 U57 ( .A(A[30]), .Y(n178) );
  INVX2 U58 ( .A(A[8]), .Y(n179) );
  INVX2 U59 ( .A(A[9]), .Y(n180) );
endmodule


module CannyEdge_DW01_add_45 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_22 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \SUMB[7][7] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] ,
         \SUMB[5][1] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] ,
         \SUMB[4][1] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , QA, QB, \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n60, n61, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign PRODUCT[1] = \ab[0][1] ;
  assign QA = TC;

  AND2X2 U2 ( .A(n41), .B(n66), .Y(n3) );
  AND2X2 U3 ( .A(n19), .B(n66), .Y(n4) );
  AND2X2 U4 ( .A(\ab[2][6] ), .B(n66), .Y(n5) );
  AND2X2 U5 ( .A(n30), .B(\SUMB[4][5] ), .Y(n6) );
  AND2X2 U6 ( .A(n28), .B(\SUMB[4][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n29), .B(\SUMB[5][2] ), .Y(n8) );
  AND2X2 U8 ( .A(n33), .B(\SUMB[2][2] ), .Y(n9) );
  AND2X2 U9 ( .A(n34), .B(\SUMB[2][3] ), .Y(n10) );
  AND2X2 U10 ( .A(n35), .B(\SUMB[2][4] ), .Y(n11) );
  AND2X2 U11 ( .A(n36), .B(\SUMB[2][5] ), .Y(n12) );
  AND2X2 U12 ( .A(n40), .B(\SUMB[6][1] ), .Y(n13) );
  AND2X2 U13 ( .A(n25), .B(\SUMB[6][3] ), .Y(n14) );
  AND2X2 U14 ( .A(n26), .B(\SUMB[6][4] ), .Y(n15) );
  AND2X2 U15 ( .A(n31), .B(\SUMB[6][5] ), .Y(n16) );
  AND2X2 U16 ( .A(\SUMB[3][1] ), .B(n39), .Y(n17) );
  AND2X2 U17 ( .A(QA), .B(QB), .Y(n18) );
  AND2X2 U18 ( .A(n3), .B(n66), .Y(n19) );
  AND2X2 U19 ( .A(\ab[0][2] ), .B(\ab[2][0] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][5] ), .B(\ab[0][7] ), .Y(n21) );
  AND2X2 U21 ( .A(n8), .B(\SUMB[6][2] ), .Y(n22) );
  AND2X2 U22 ( .A(n11), .B(\SUMB[3][4] ), .Y(n23) );
  AND2X2 U23 ( .A(n23), .B(\SUMB[4][4] ), .Y(n24) );
  AND2X2 U24 ( .A(n7), .B(\SUMB[5][3] ), .Y(n25) );
  AND2X2 U25 ( .A(n24), .B(\SUMB[5][4] ), .Y(n26) );
  AND2X2 U26 ( .A(n9), .B(\SUMB[3][2] ), .Y(n27) );
  AND2X2 U27 ( .A(n10), .B(\SUMB[3][3] ), .Y(n28) );
  AND2X2 U28 ( .A(n27), .B(\SUMB[4][2] ), .Y(n29) );
  AND2X2 U29 ( .A(n12), .B(\SUMB[3][5] ), .Y(n30) );
  AND2X2 U30 ( .A(n6), .B(\SUMB[5][5] ), .Y(n31) );
  AND2X2 U31 ( .A(n21), .B(\SUMB[2][6] ), .Y(n32) );
  AND2X2 U32 ( .A(\ab[2][1] ), .B(\ab[0][3] ), .Y(n33) );
  AND2X2 U33 ( .A(\ab[2][2] ), .B(\ab[0][4] ), .Y(n34) );
  AND2X2 U34 ( .A(\ab[2][3] ), .B(\ab[0][5] ), .Y(n35) );
  AND2X2 U35 ( .A(\ab[2][4] ), .B(\ab[0][6] ), .Y(n36) );
  AND2X2 U36 ( .A(\SUMB[7][1] ), .B(n13), .Y(n37) );
  AND2X2 U37 ( .A(\SUMB[4][1] ), .B(n17), .Y(n38) );
  AND2X2 U38 ( .A(\SUMB[2][1] ), .B(n20), .Y(n39) );
  AND2X2 U39 ( .A(\SUMB[5][1] ), .B(n38), .Y(n40) );
  AND2X2 U40 ( .A(n32), .B(n5), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[7][0] ), .B(n66), .Y(n42) );
  AND2X2 U42 ( .A(n66), .B(n4), .Y(n43) );
  AND2X2 U43 ( .A(\SUMB[7][3] ), .B(n14), .Y(n44) );
  AND2X2 U44 ( .A(\SUMB[7][2] ), .B(n22), .Y(n45) );
  AND2X2 U45 ( .A(\SUMB[7][4] ), .B(n15), .Y(n46) );
  AND2X2 U46 ( .A(\SUMB[7][5] ), .B(n16), .Y(n47) );
  XOR2X1 U47 ( .A(\SUMB[7][1] ), .B(n13), .Y(\A1[6] ) );
  XOR2X1 U48 ( .A(\SUMB[7][2] ), .B(n22), .Y(\A1[7] ) );
  XOR2X1 U49 ( .A(\SUMB[7][3] ), .B(n14), .Y(\A1[8] ) );
  XOR2X1 U50 ( .A(\SUMB[7][4] ), .B(n15), .Y(\A1[9] ) );
  XOR2X1 U51 ( .A(\SUMB[7][5] ), .B(n16), .Y(\A1[10] ) );
  XOR2X1 U52 ( .A(n66), .B(n4), .Y(\A1[11] ) );
  XOR2X1 U53 ( .A(n18), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U54 ( .A(\SUMB[7][0] ), .B(n66), .Y(\A1[5] ) );
  XOR2X1 U55 ( .A(\SUMB[2][1] ), .B(n20), .Y(\A1[1] ) );
  XOR2X1 U56 ( .A(\SUMB[2][2] ), .B(n33), .Y(\SUMB[3][1] ) );
  XOR2X1 U57 ( .A(\SUMB[2][3] ), .B(n34), .Y(\SUMB[3][2] ) );
  XOR2X1 U58 ( .A(\SUMB[2][4] ), .B(n35), .Y(\SUMB[3][3] ) );
  XOR2X1 U59 ( .A(\SUMB[2][5] ), .B(n36), .Y(\SUMB[3][4] ) );
  XOR2X1 U60 ( .A(\SUMB[2][6] ), .B(n21), .Y(\SUMB[3][5] ) );
  XOR2X1 U61 ( .A(\SUMB[3][1] ), .B(n39), .Y(\A1[2] ) );
  XOR2X1 U62 ( .A(\SUMB[3][2] ), .B(n9), .Y(\SUMB[4][1] ) );
  XOR2X1 U63 ( .A(\SUMB[3][3] ), .B(n10), .Y(\SUMB[4][2] ) );
  XOR2X1 U64 ( .A(\SUMB[3][4] ), .B(n11), .Y(\SUMB[4][3] ) );
  XOR2X1 U65 ( .A(\SUMB[3][5] ), .B(n12), .Y(\SUMB[4][4] ) );
  XOR2X1 U66 ( .A(n5), .B(n32), .Y(\SUMB[4][5] ) );
  XOR2X1 U67 ( .A(\SUMB[4][1] ), .B(n17), .Y(\A1[3] ) );
  XOR2X1 U68 ( .A(\SUMB[4][2] ), .B(n27), .Y(\SUMB[5][1] ) );
  XOR2X1 U69 ( .A(\SUMB[4][3] ), .B(n28), .Y(\SUMB[5][2] ) );
  XOR2X1 U70 ( .A(\SUMB[4][4] ), .B(n23), .Y(\SUMB[5][3] ) );
  XOR2X1 U71 ( .A(\SUMB[4][5] ), .B(n30), .Y(\SUMB[5][4] ) );
  XOR2X1 U72 ( .A(n66), .B(n41), .Y(\SUMB[5][5] ) );
  XOR2X1 U73 ( .A(\SUMB[5][1] ), .B(n38), .Y(\A1[4] ) );
  XOR2X1 U74 ( .A(\SUMB[5][2] ), .B(n29), .Y(\SUMB[6][1] ) );
  XOR2X1 U75 ( .A(\SUMB[5][3] ), .B(n7), .Y(\SUMB[6][2] ) );
  XOR2X1 U76 ( .A(\SUMB[5][4] ), .B(n24), .Y(\SUMB[6][3] ) );
  XOR2X1 U77 ( .A(\SUMB[5][5] ), .B(n6), .Y(\SUMB[6][4] ) );
  XOR2X1 U78 ( .A(n66), .B(n3), .Y(\SUMB[6][5] ) );
  XOR2X1 U79 ( .A(\SUMB[6][1] ), .B(n40), .Y(\SUMB[7][0] ) );
  XOR2X1 U80 ( .A(\SUMB[6][2] ), .B(n8), .Y(\SUMB[7][1] ) );
  XOR2X1 U81 ( .A(\SUMB[6][3] ), .B(n25), .Y(\SUMB[7][2] ) );
  XOR2X1 U82 ( .A(\SUMB[6][4] ), .B(n26), .Y(\SUMB[7][3] ) );
  XOR2X1 U83 ( .A(\SUMB[6][5] ), .B(n31), .Y(\SUMB[7][4] ) );
  XOR2X1 U84 ( .A(n66), .B(n19), .Y(\SUMB[7][5] ) );
  XOR2X1 U85 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  XOR2X1 U86 ( .A(\ab[0][2] ), .B(\ab[2][0] ), .Y(\A1[0] ) );
  XOR2X1 U87 ( .A(\ab[0][3] ), .B(\ab[2][1] ), .Y(\SUMB[2][1] ) );
  XOR2X1 U88 ( .A(\ab[0][4] ), .B(\ab[2][2] ), .Y(\SUMB[2][2] ) );
  XOR2X1 U89 ( .A(\ab[0][5] ), .B(\ab[2][3] ), .Y(\SUMB[2][3] ) );
  XOR2X1 U90 ( .A(\ab[0][6] ), .B(\ab[2][4] ), .Y(\SUMB[2][4] ) );
  XOR2X1 U91 ( .A(\ab[0][7] ), .B(\ab[2][5] ), .Y(\SUMB[2][5] ) );
  XOR2X1 U92 ( .A(n66), .B(\ab[2][6] ), .Y(\SUMB[2][6] ) );
  NOR2X1 U104 ( .A(n65), .B(n72), .Y(\ab[2][6] ) );
  NOR2X1 U105 ( .A(n65), .B(n71), .Y(\ab[2][5] ) );
  NOR2X1 U106 ( .A(n65), .B(n70), .Y(\ab[2][4] ) );
  NOR2X1 U107 ( .A(n65), .B(n69), .Y(\ab[2][3] ) );
  NOR2X1 U108 ( .A(n65), .B(n68), .Y(\ab[2][2] ) );
  NOR2X1 U109 ( .A(n65), .B(n67), .Y(\ab[2][1] ) );
  NOR2X1 U110 ( .A(n65), .B(n74), .Y(\ab[2][0] ) );
  MUX2X1 U111 ( .B(n60), .A(n61), .S(A[0]), .Y(\ab[0][7] ) );
  NAND2X1 U112 ( .A(B[7]), .B(n65), .Y(n61) );
  NOR2X1 U113 ( .A(n72), .B(n73), .Y(\ab[0][6] ) );
  NOR2X1 U114 ( .A(n71), .B(n73), .Y(\ab[0][5] ) );
  NOR2X1 U115 ( .A(n70), .B(n73), .Y(\ab[0][4] ) );
  NOR2X1 U116 ( .A(n69), .B(n73), .Y(\ab[0][3] ) );
  NOR2X1 U117 ( .A(n68), .B(n73), .Y(\ab[0][2] ) );
  NOR2X1 U118 ( .A(n67), .B(n73), .Y(\ab[0][1] ) );
  NAND2X1 U119 ( .A(QA), .B(B[7]), .Y(n60) );
  NOR2X1 U120 ( .A(B[7]), .B(n65), .Y(QB) );
  NOR2X1 U121 ( .A(n74), .B(n73), .Y(PRODUCT[0]) );
  CannyEdge_DW01_add_45 FS_1 ( .A({\A1[13] , \SUMB[7][7] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({1'b0, n43, n47, n46, n44, n45, n37, n42, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U96 ( .A(QA), .Y(n65) );
  INVX2 U97 ( .A(n60), .Y(n66) );
  INVX2 U98 ( .A(B[1]), .Y(n67) );
  INVX2 U99 ( .A(B[2]), .Y(n68) );
  INVX2 U100 ( .A(B[3]), .Y(n69) );
  INVX2 U101 ( .A(B[4]), .Y(n70) );
  INVX2 U102 ( .A(B[5]), .Y(n71) );
  INVX2 U103 ( .A(B[6]), .Y(n72) );
  INVX2 U122 ( .A(A[0]), .Y(n73) );
  INVX2 U123 ( .A(B[0]), .Y(n74) );
endmodule


module CannyEdge_DW01_add_47 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40;
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X1 U11 ( .A(n10), .B(n11), .Y(SUM[9]) );
  NOR2X1 U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n14), .B(n37), .Y(SUM[8]) );
  NAND2X1 U14 ( .A(n36), .B(n15), .Y(n14) );
  XOR2X1 U15 ( .A(n17), .B(n18), .Y(SUM[7]) );
  XOR2X1 U16 ( .A(n38), .B(B[7]), .Y(n18) );
  OAI21X1 U17 ( .A(B[6]), .B(A[6]), .C(n17), .Y(n19) );
  XOR2X1 U18 ( .A(n20), .B(n21), .Y(SUM[12]) );
  XOR2X1 U19 ( .A(B[12]), .B(A[12]), .Y(n21) );
  OAI21X1 U20 ( .A(n22), .B(n33), .C(n23), .Y(n20) );
  XOR2X1 U21 ( .A(n24), .B(n25), .Y(SUM[11]) );
  NOR2X1 U22 ( .A(n32), .B(n22), .Y(n25) );
  NOR2X1 U23 ( .A(B[11]), .B(A[11]), .Y(n22) );
  NAND2X1 U24 ( .A(B[11]), .B(A[11]), .Y(n23) );
  OAI21X1 U25 ( .A(n26), .B(n27), .C(n28), .Y(n24) );
  XOR2X1 U26 ( .A(n29), .B(n27), .Y(SUM[10]) );
  AOI21X1 U27 ( .A(n10), .B(n35), .C(n12), .Y(n27) );
  AND2X1 U28 ( .A(B[9]), .B(A[9]), .Y(n12) );
  NOR2X1 U29 ( .A(B[9]), .B(A[9]), .Y(n13) );
  OAI21X1 U30 ( .A(n37), .B(n16), .C(n15), .Y(n10) );
  NAND2X1 U31 ( .A(B[8]), .B(A[8]), .Y(n15) );
  NOR2X1 U32 ( .A(B[8]), .B(A[8]), .Y(n16) );
  OAI21X1 U33 ( .A(n17), .B(n38), .C(n31), .Y(n30) );
  OAI21X1 U34 ( .A(n40), .B(A[7]), .C(B[7]), .Y(n31) );
  NAND2X1 U35 ( .A(B[6]), .B(A[6]), .Y(n17) );
  NAND2X1 U36 ( .A(n34), .B(n28), .Y(n29) );
  NAND2X1 U37 ( .A(B[10]), .B(A[10]), .Y(n28) );
  NOR2X1 U38 ( .A(B[10]), .B(A[10]), .Y(n26) );
  INVX2 U2 ( .A(n23), .Y(n32) );
  INVX2 U3 ( .A(n24), .Y(n33) );
  INVX2 U4 ( .A(n26), .Y(n34) );
  INVX2 U5 ( .A(n13), .Y(n35) );
  INVX2 U6 ( .A(n16), .Y(n36) );
  INVX2 U7 ( .A(n30), .Y(n37) );
  INVX2 U8 ( .A(A[7]), .Y(n38) );
  INVX2 U9 ( .A(n19), .Y(SUM[6]) );
  INVX2 U10 ( .A(n17), .Y(n40) );
endmodule


module CannyEdge_DW02_mult_23 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] ,
         \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] ,
         \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , QA, QB,
         \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] ,
         \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n57, n58, n61, n62;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign PRODUCT[0] = \ab[2][0] ;
  assign QA = TC;

  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n23), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n22), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n21), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n20), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n19), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n18), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  FAX1 S3_2_6 ( .A(\ab[2][6] ), .B(n24), .C(\ab[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  AND2X2 U2 ( .A(\SUMB[7][7] ), .B(n5), .Y(n3) );
  AND2X2 U3 ( .A(n28), .B(n62), .Y(n4) );
  AND2X2 U4 ( .A(n27), .B(n62), .Y(n5) );
  AND2X2 U5 ( .A(n43), .B(\SUMB[3][2] ), .Y(n6) );
  AND2X2 U6 ( .A(n44), .B(\SUMB[3][3] ), .Y(n7) );
  AND2X2 U7 ( .A(n45), .B(\SUMB[3][4] ), .Y(n8) );
  AND2X2 U8 ( .A(n46), .B(\SUMB[3][5] ), .Y(n9) );
  AND2X2 U9 ( .A(n47), .B(\SUMB[3][6] ), .Y(n10) );
  AND2X2 U10 ( .A(n42), .B(\SUMB[6][1] ), .Y(n11) );
  AND2X2 U11 ( .A(n34), .B(\SUMB[6][2] ), .Y(n12) );
  AND2X2 U12 ( .A(n35), .B(\SUMB[6][3] ), .Y(n13) );
  AND2X2 U13 ( .A(n36), .B(\SUMB[6][4] ), .Y(n14) );
  AND2X2 U14 ( .A(n37), .B(\SUMB[6][5] ), .Y(n15) );
  AND2X2 U15 ( .A(n39), .B(\SUMB[6][6] ), .Y(n16) );
  AND2X2 U16 ( .A(\SUMB[4][1] ), .B(n41), .Y(n17) );
  AND2X2 U17 ( .A(\ab[2][6] ), .B(\ab[1][5] ), .Y(n18) );
  AND2X2 U18 ( .A(\ab[2][5] ), .B(\ab[1][4] ), .Y(n19) );
  AND2X2 U19 ( .A(\ab[2][4] ), .B(\ab[1][3] ), .Y(n20) );
  AND2X2 U20 ( .A(\ab[2][3] ), .B(\ab[1][2] ), .Y(n21) );
  AND2X2 U21 ( .A(\ab[2][2] ), .B(\ab[1][1] ), .Y(n22) );
  AND2X2 U22 ( .A(\ab[2][1] ), .B(\ab[1][0] ), .Y(n23) );
  AND2X2 U23 ( .A(\ab[2][7] ), .B(\ab[1][6] ), .Y(n24) );
  AND2X2 U24 ( .A(QA), .B(QB), .Y(n25) );
  AND2X2 U25 ( .A(n4), .B(n62), .Y(n26) );
  AND2X2 U26 ( .A(n26), .B(n62), .Y(n27) );
  AND2X2 U27 ( .A(\CARRYB[2][6] ), .B(\ab[2][7] ), .Y(n28) );
  AND2X2 U28 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(n29) );
  AND2X2 U29 ( .A(n6), .B(\SUMB[4][2] ), .Y(n30) );
  AND2X2 U30 ( .A(n7), .B(\SUMB[4][3] ), .Y(n31) );
  AND2X2 U31 ( .A(n8), .B(\SUMB[4][4] ), .Y(n32) );
  AND2X2 U32 ( .A(n9), .B(\SUMB[4][5] ), .Y(n33) );
  AND2X2 U33 ( .A(n30), .B(\SUMB[5][2] ), .Y(n34) );
  AND2X2 U34 ( .A(n31), .B(\SUMB[5][3] ), .Y(n35) );
  AND2X2 U35 ( .A(n32), .B(\SUMB[5][4] ), .Y(n36) );
  AND2X2 U36 ( .A(n33), .B(\SUMB[5][5] ), .Y(n37) );
  AND2X2 U37 ( .A(n10), .B(\SUMB[4][6] ), .Y(n38) );
  AND2X2 U38 ( .A(n38), .B(\SUMB[5][6] ), .Y(n39) );
  AND2X2 U39 ( .A(\SUMB[7][1] ), .B(n11), .Y(n40) );
  AND2X2 U40 ( .A(\SUMB[3][1] ), .B(n29), .Y(n41) );
  AND2X2 U41 ( .A(\SUMB[5][1] ), .B(n17), .Y(n42) );
  AND2X2 U42 ( .A(\CARRYB[2][1] ), .B(\SUMB[2][2] ), .Y(n43) );
  AND2X2 U43 ( .A(\CARRYB[2][2] ), .B(\SUMB[2][3] ), .Y(n44) );
  AND2X2 U44 ( .A(\CARRYB[2][3] ), .B(\SUMB[2][4] ), .Y(n45) );
  AND2X2 U45 ( .A(\CARRYB[2][4] ), .B(\SUMB[2][5] ), .Y(n46) );
  AND2X2 U46 ( .A(\CARRYB[2][5] ), .B(\SUMB[2][6] ), .Y(n47) );
  AND2X2 U47 ( .A(\SUMB[7][0] ), .B(n62), .Y(n48) );
  AND2X2 U48 ( .A(\SUMB[7][6] ), .B(n16), .Y(n49) );
  AND2X2 U49 ( .A(\SUMB[7][3] ), .B(n13), .Y(n50) );
  AND2X2 U50 ( .A(\SUMB[7][5] ), .B(n15), .Y(n51) );
  AND2X2 U51 ( .A(\SUMB[7][2] ), .B(n12), .Y(n52) );
  AND2X2 U52 ( .A(\SUMB[7][4] ), .B(n14), .Y(n53) );
  XOR2X1 U53 ( .A(\SUMB[7][1] ), .B(n11), .Y(\A1[6] ) );
  XOR2X1 U54 ( .A(\SUMB[7][2] ), .B(n12), .Y(\A1[7] ) );
  XOR2X1 U55 ( .A(\SUMB[7][3] ), .B(n13), .Y(\A1[8] ) );
  XOR2X1 U56 ( .A(\SUMB[7][4] ), .B(n14), .Y(\A1[9] ) );
  XOR2X1 U57 ( .A(\SUMB[7][5] ), .B(n15), .Y(\A1[10] ) );
  XOR2X1 U58 ( .A(\SUMB[7][6] ), .B(n16), .Y(\A1[11] ) );
  XOR2X1 U59 ( .A(\SUMB[7][7] ), .B(n5), .Y(\A1[12] ) );
  XOR2X1 U60 ( .A(n25), .B(QA), .Y(\A1[13] ) );
  XOR2X1 U61 ( .A(\ab[1][0] ), .B(\ab[2][1] ), .Y(PRODUCT[1]) );
  XOR2X1 U62 ( .A(\ab[1][1] ), .B(\ab[2][2] ), .Y(\SUMB[1][1] ) );
  XOR2X1 U63 ( .A(\ab[1][2] ), .B(\ab[2][3] ), .Y(\SUMB[1][2] ) );
  XOR2X1 U64 ( .A(\ab[1][3] ), .B(\ab[2][4] ), .Y(\SUMB[1][3] ) );
  XOR2X1 U65 ( .A(\ab[1][4] ), .B(\ab[2][5] ), .Y(\SUMB[1][4] ) );
  XOR2X1 U66 ( .A(\ab[1][5] ), .B(\ab[2][6] ), .Y(\SUMB[1][5] ) );
  XOR2X1 U67 ( .A(\ab[1][6] ), .B(\ab[2][7] ), .Y(\SUMB[1][6] ) );
  XOR2X1 U68 ( .A(\SUMB[7][0] ), .B(n62), .Y(\A1[5] ) );
  XOR2X1 U69 ( .A(\SUMB[2][1] ), .B(\CARRYB[2][0] ), .Y(\A1[1] ) );
  XOR2X1 U70 ( .A(\SUMB[2][2] ), .B(\CARRYB[2][1] ), .Y(\SUMB[3][1] ) );
  XOR2X1 U71 ( .A(\SUMB[2][3] ), .B(\CARRYB[2][2] ), .Y(\SUMB[3][2] ) );
  XOR2X1 U72 ( .A(\SUMB[2][4] ), .B(\CARRYB[2][3] ), .Y(\SUMB[3][3] ) );
  XOR2X1 U73 ( .A(\SUMB[2][5] ), .B(\CARRYB[2][4] ), .Y(\SUMB[3][4] ) );
  XOR2X1 U74 ( .A(\SUMB[2][6] ), .B(\CARRYB[2][5] ), .Y(\SUMB[3][5] ) );
  XOR2X1 U75 ( .A(\ab[2][7] ), .B(\CARRYB[2][6] ), .Y(\SUMB[3][6] ) );
  XOR2X1 U76 ( .A(\SUMB[3][1] ), .B(n29), .Y(\A1[2] ) );
  XOR2X1 U77 ( .A(\SUMB[3][2] ), .B(n43), .Y(\SUMB[4][1] ) );
  XOR2X1 U78 ( .A(\SUMB[3][3] ), .B(n44), .Y(\SUMB[4][2] ) );
  XOR2X1 U79 ( .A(\SUMB[3][4] ), .B(n45), .Y(\SUMB[4][3] ) );
  XOR2X1 U80 ( .A(\SUMB[3][5] ), .B(n46), .Y(\SUMB[4][4] ) );
  XOR2X1 U81 ( .A(\SUMB[3][6] ), .B(n47), .Y(\SUMB[4][5] ) );
  XOR2X1 U82 ( .A(n62), .B(n28), .Y(\SUMB[4][6] ) );
  XOR2X1 U83 ( .A(\SUMB[4][1] ), .B(n41), .Y(\A1[3] ) );
  XOR2X1 U84 ( .A(\SUMB[4][2] ), .B(n6), .Y(\SUMB[5][1] ) );
  XOR2X1 U85 ( .A(\SUMB[4][3] ), .B(n7), .Y(\SUMB[5][2] ) );
  XOR2X1 U86 ( .A(\SUMB[4][4] ), .B(n8), .Y(\SUMB[5][3] ) );
  XOR2X1 U87 ( .A(\SUMB[4][5] ), .B(n9), .Y(\SUMB[5][4] ) );
  XOR2X1 U88 ( .A(\SUMB[4][6] ), .B(n10), .Y(\SUMB[5][5] ) );
  XOR2X1 U89 ( .A(n62), .B(n4), .Y(\SUMB[5][6] ) );
  XOR2X1 U90 ( .A(\SUMB[5][1] ), .B(n17), .Y(\A1[4] ) );
  XOR2X1 U91 ( .A(\SUMB[5][2] ), .B(n30), .Y(\SUMB[6][1] ) );
  XOR2X1 U92 ( .A(\SUMB[5][3] ), .B(n31), .Y(\SUMB[6][2] ) );
  XOR2X1 U93 ( .A(\SUMB[5][4] ), .B(n32), .Y(\SUMB[6][3] ) );
  XOR2X1 U94 ( .A(\SUMB[5][5] ), .B(n33), .Y(\SUMB[6][4] ) );
  XOR2X1 U95 ( .A(\SUMB[5][6] ), .B(n38), .Y(\SUMB[6][5] ) );
  XOR2X1 U96 ( .A(n62), .B(n26), .Y(\SUMB[6][6] ) );
  XOR2X1 U97 ( .A(\SUMB[6][1] ), .B(n42), .Y(\SUMB[7][0] ) );
  XOR2X1 U98 ( .A(\SUMB[6][2] ), .B(n34), .Y(\SUMB[7][1] ) );
  XOR2X1 U99 ( .A(\SUMB[6][3] ), .B(n35), .Y(\SUMB[7][2] ) );
  XOR2X1 U100 ( .A(\SUMB[6][4] ), .B(n36), .Y(\SUMB[7][3] ) );
  XOR2X1 U101 ( .A(\SUMB[6][5] ), .B(n37), .Y(\SUMB[7][4] ) );
  XOR2X1 U102 ( .A(\SUMB[6][6] ), .B(n39), .Y(\SUMB[7][5] ) );
  XOR2X1 U103 ( .A(n62), .B(n27), .Y(\SUMB[7][6] ) );
  XOR2X1 U104 ( .A(QB), .B(QA), .Y(\SUMB[7][7] ) );
  MUX2X1 U107 ( .B(n57), .A(n58), .S(A[1]), .Y(\ab[1][7] ) );
  AND2X1 U108 ( .A(B[6]), .B(A[1]), .Y(\ab[1][6] ) );
  AND2X1 U109 ( .A(B[5]), .B(A[1]), .Y(\ab[1][5] ) );
  AND2X1 U110 ( .A(B[4]), .B(A[1]), .Y(\ab[1][4] ) );
  AND2X1 U111 ( .A(B[3]), .B(A[1]), .Y(\ab[1][3] ) );
  AND2X1 U112 ( .A(B[2]), .B(A[1]), .Y(\ab[1][2] ) );
  AND2X1 U113 ( .A(B[1]), .B(A[1]), .Y(\ab[1][1] ) );
  AND2X1 U114 ( .A(B[0]), .B(A[1]), .Y(\ab[1][0] ) );
  MUX2X1 U115 ( .B(n57), .A(n58), .S(A[2]), .Y(\ab[2][7] ) );
  NAND2X1 U116 ( .A(B[7]), .B(n61), .Y(n58) );
  AND2X1 U117 ( .A(B[6]), .B(A[2]), .Y(\ab[2][6] ) );
  AND2X1 U118 ( .A(B[5]), .B(A[2]), .Y(\ab[2][5] ) );
  AND2X1 U119 ( .A(B[4]), .B(A[2]), .Y(\ab[2][4] ) );
  AND2X1 U120 ( .A(B[3]), .B(A[2]), .Y(\ab[2][3] ) );
  AND2X1 U121 ( .A(B[2]), .B(A[2]), .Y(\ab[2][2] ) );
  AND2X1 U122 ( .A(B[1]), .B(A[2]), .Y(\ab[2][1] ) );
  NAND2X1 U123 ( .A(QA), .B(B[7]), .Y(n57) );
  NOR2X1 U124 ( .A(B[7]), .B(n61), .Y(QB) );
  AND2X1 U125 ( .A(B[0]), .B(A[2]), .Y(\ab[2][0] ) );
  CannyEdge_DW01_add_47 FS_1 ( .A({\A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({n3, n49, n51, n53, n50, n52, n40, n48, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, PRODUCT[14:2]}) );
  INVX2 U126 ( .A(QA), .Y(n61) );
  INVX2 U127 ( .A(n57), .Y(n62) );
endmodule


module CannyEdge_DW01_cmp2_6 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188;

  MUX2X1 U63 ( .B(n63), .A(n64), .S(B[31]), .Y(LT_LE) );
  MUX2X1 U64 ( .B(n160), .A(n65), .S(A[31]), .Y(n64) );
  NOR2X1 U65 ( .A(n66), .B(n186), .Y(n65) );
  MUX2X1 U66 ( .B(n67), .A(TC), .S(A[31]), .Y(n63) );
  NAND2X1 U67 ( .A(n66), .B(n186), .Y(n67) );
  AOI21X1 U68 ( .A(n134), .B(B[29]), .C(n127), .Y(n66) );
  OAI21X1 U69 ( .A(B[29]), .B(n134), .C(n69), .Y(n68) );
  AOI21X1 U70 ( .A(A[28]), .B(n185), .C(n70), .Y(n69) );
  AOI21X1 U71 ( .A(B[28]), .B(n135), .C(n71), .Y(n70) );
  OAI21X1 U72 ( .A(A[27]), .B(n184), .C(n72), .Y(n71) );
  OAI21X1 U73 ( .A(B[27]), .B(n136), .C(n73), .Y(n72) );
  AOI21X1 U74 ( .A(A[26]), .B(n183), .C(n74), .Y(n73) );
  AOI21X1 U75 ( .A(B[26]), .B(n137), .C(n75), .Y(n74) );
  OAI21X1 U76 ( .A(A[25]), .B(n182), .C(n76), .Y(n75) );
  OAI21X1 U77 ( .A(B[25]), .B(n138), .C(n77), .Y(n76) );
  AOI21X1 U78 ( .A(A[24]), .B(n181), .C(n78), .Y(n77) );
  AOI21X1 U79 ( .A(B[24]), .B(n139), .C(n79), .Y(n78) );
  OAI21X1 U80 ( .A(A[23]), .B(n180), .C(n80), .Y(n79) );
  OAI21X1 U81 ( .A(B[23]), .B(n140), .C(n81), .Y(n80) );
  AOI21X1 U82 ( .A(A[22]), .B(n179), .C(n82), .Y(n81) );
  AOI21X1 U83 ( .A(B[22]), .B(n141), .C(n83), .Y(n82) );
  OAI21X1 U84 ( .A(A[21]), .B(n178), .C(n84), .Y(n83) );
  OAI21X1 U85 ( .A(B[21]), .B(n142), .C(n85), .Y(n84) );
  AOI21X1 U86 ( .A(A[20]), .B(n177), .C(n86), .Y(n85) );
  AOI21X1 U87 ( .A(B[20]), .B(n143), .C(n87), .Y(n86) );
  OAI21X1 U88 ( .A(A[19]), .B(n176), .C(n88), .Y(n87) );
  OAI21X1 U89 ( .A(B[19]), .B(n144), .C(n89), .Y(n88) );
  AOI21X1 U90 ( .A(A[18]), .B(n175), .C(n90), .Y(n89) );
  AOI21X1 U91 ( .A(B[18]), .B(n145), .C(n91), .Y(n90) );
  OAI21X1 U92 ( .A(A[17]), .B(n174), .C(n92), .Y(n91) );
  OAI21X1 U93 ( .A(B[17]), .B(n146), .C(n93), .Y(n92) );
  AOI21X1 U94 ( .A(A[16]), .B(n173), .C(n94), .Y(n93) );
  AOI21X1 U95 ( .A(B[16]), .B(n147), .C(n95), .Y(n94) );
  OAI21X1 U96 ( .A(A[15]), .B(n172), .C(n96), .Y(n95) );
  OAI21X1 U97 ( .A(B[15]), .B(n148), .C(n97), .Y(n96) );
  AOI21X1 U98 ( .A(A[14]), .B(n171), .C(n98), .Y(n97) );
  AOI21X1 U99 ( .A(B[14]), .B(n149), .C(n99), .Y(n98) );
  OAI21X1 U100 ( .A(A[13]), .B(n170), .C(n100), .Y(n99) );
  OAI21X1 U101 ( .A(B[13]), .B(n150), .C(n101), .Y(n100) );
  AOI21X1 U102 ( .A(A[12]), .B(n169), .C(n102), .Y(n101) );
  AOI21X1 U103 ( .A(B[12]), .B(n151), .C(n103), .Y(n102) );
  OAI21X1 U104 ( .A(A[11]), .B(n168), .C(n104), .Y(n103) );
  OAI21X1 U105 ( .A(B[11]), .B(n152), .C(n105), .Y(n104) );
  AOI21X1 U106 ( .A(A[10]), .B(n167), .C(n106), .Y(n105) );
  AOI21X1 U107 ( .A(B[10]), .B(n153), .C(n107), .Y(n106) );
  OAI21X1 U108 ( .A(A[9]), .B(n188), .C(n108), .Y(n107) );
  OAI21X1 U109 ( .A(B[9]), .B(n154), .C(n109), .Y(n108) );
  AOI21X1 U110 ( .A(A[8]), .B(n187), .C(n110), .Y(n109) );
  AOI21X1 U111 ( .A(B[8]), .B(n155), .C(n111), .Y(n110) );
  OAI21X1 U112 ( .A(A[7]), .B(n161), .C(n112), .Y(n111) );
  OAI21X1 U113 ( .A(B[7]), .B(n156), .C(n113), .Y(n112) );
  AOI21X1 U114 ( .A(A[6]), .B(n162), .C(n114), .Y(n113) );
  AOI21X1 U115 ( .A(B[6]), .B(n157), .C(n115), .Y(n114) );
  OAI21X1 U116 ( .A(A[5]), .B(n163), .C(n116), .Y(n115) );
  OAI21X1 U117 ( .A(B[5]), .B(n158), .C(n117), .Y(n116) );
  AOI21X1 U118 ( .A(A[4]), .B(n164), .C(n118), .Y(n117) );
  AOI21X1 U119 ( .A(B[4]), .B(n159), .C(n119), .Y(n118) );
  OAI21X1 U120 ( .A(A[3]), .B(n133), .C(n120), .Y(n119) );
  OAI21X1 U121 ( .A(B[3]), .B(n131), .C(n121), .Y(n120) );
  AOI21X1 U122 ( .A(A[2]), .B(n165), .C(n122), .Y(n121) );
  AOI21X1 U123 ( .A(B[2]), .B(n130), .C(n123), .Y(n122) );
  OAI21X1 U124 ( .A(A[1]), .B(n132), .C(n124), .Y(n123) );
  OAI21X1 U125 ( .A(B[1]), .B(n129), .C(n125), .Y(n124) );
  AOI21X1 U126 ( .A(A[0]), .B(n166), .C(n126), .Y(n125) );
  AOI21X1 U127 ( .A(B[0]), .B(n128), .C(LEQ), .Y(n126) );
  INVX2 U1 ( .A(n68), .Y(n127) );
  INVX2 U2 ( .A(A[0]), .Y(n128) );
  INVX2 U3 ( .A(A[1]), .Y(n129) );
  INVX2 U4 ( .A(A[2]), .Y(n130) );
  INVX2 U5 ( .A(A[3]), .Y(n131) );
  INVX2 U6 ( .A(B[1]), .Y(n132) );
  INVX2 U7 ( .A(B[3]), .Y(n133) );
  INVX2 U8 ( .A(A[29]), .Y(n134) );
  INVX2 U9 ( .A(A[28]), .Y(n135) );
  INVX2 U10 ( .A(A[27]), .Y(n136) );
  INVX2 U11 ( .A(A[26]), .Y(n137) );
  INVX2 U12 ( .A(A[25]), .Y(n138) );
  INVX2 U13 ( .A(A[24]), .Y(n139) );
  INVX2 U14 ( .A(A[23]), .Y(n140) );
  INVX2 U15 ( .A(A[22]), .Y(n141) );
  INVX2 U16 ( .A(A[21]), .Y(n142) );
  INVX2 U17 ( .A(A[20]), .Y(n143) );
  INVX2 U18 ( .A(A[19]), .Y(n144) );
  INVX2 U19 ( .A(A[18]), .Y(n145) );
  INVX2 U20 ( .A(A[17]), .Y(n146) );
  INVX2 U21 ( .A(A[16]), .Y(n147) );
  INVX2 U22 ( .A(A[15]), .Y(n148) );
  INVX2 U23 ( .A(A[14]), .Y(n149) );
  INVX2 U24 ( .A(A[13]), .Y(n150) );
  INVX2 U25 ( .A(A[12]), .Y(n151) );
  INVX2 U26 ( .A(A[11]), .Y(n152) );
  INVX2 U27 ( .A(A[10]), .Y(n153) );
  INVX2 U28 ( .A(A[9]), .Y(n154) );
  INVX2 U29 ( .A(A[8]), .Y(n155) );
  INVX2 U30 ( .A(A[7]), .Y(n156) );
  INVX2 U31 ( .A(A[6]), .Y(n157) );
  INVX2 U32 ( .A(A[5]), .Y(n158) );
  INVX2 U33 ( .A(A[4]), .Y(n159) );
  INVX2 U34 ( .A(TC), .Y(n160) );
  INVX2 U35 ( .A(B[7]), .Y(n161) );
  INVX2 U36 ( .A(B[6]), .Y(n162) );
  INVX2 U37 ( .A(B[5]), .Y(n163) );
  INVX2 U38 ( .A(B[4]), .Y(n164) );
  INVX2 U39 ( .A(B[2]), .Y(n165) );
  INVX2 U40 ( .A(B[0]), .Y(n166) );
  INVX2 U41 ( .A(B[10]), .Y(n167) );
  INVX2 U42 ( .A(B[11]), .Y(n168) );
  INVX2 U43 ( .A(B[12]), .Y(n169) );
  INVX2 U44 ( .A(B[13]), .Y(n170) );
  INVX2 U45 ( .A(B[14]), .Y(n171) );
  INVX2 U46 ( .A(B[15]), .Y(n172) );
  INVX2 U47 ( .A(B[16]), .Y(n173) );
  INVX2 U48 ( .A(B[17]), .Y(n174) );
  INVX2 U49 ( .A(B[18]), .Y(n175) );
  INVX2 U50 ( .A(B[19]), .Y(n176) );
  INVX2 U51 ( .A(B[20]), .Y(n177) );
  INVX2 U52 ( .A(B[21]), .Y(n178) );
  INVX2 U53 ( .A(B[22]), .Y(n179) );
  INVX2 U54 ( .A(B[23]), .Y(n180) );
  INVX2 U55 ( .A(B[24]), .Y(n181) );
  INVX2 U56 ( .A(B[25]), .Y(n182) );
  INVX2 U57 ( .A(B[26]), .Y(n183) );
  INVX2 U58 ( .A(B[27]), .Y(n184) );
  INVX2 U59 ( .A(B[28]), .Y(n185) );
  INVX2 U60 ( .A(B[30]), .Y(n186) );
  INVX2 U61 ( .A(B[8]), .Y(n187) );
  INVX2 U62 ( .A(B[9]), .Y(n188) );
endmodule


module CannyEdge_DW01_addsub_16 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [32:0] carry;
  wire   [31:0] B_AS;
  assign carry[0] = ADD_SUB;

  FAX1 U1_7 ( .A(A[7]), .B(B_AS[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7])
         );
  FAX1 U1_6 ( .A(A[6]), .B(B_AS[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6])
         );
  FAX1 U1_5 ( .A(A[5]), .B(B_AS[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5])
         );
  FAX1 U1_4 ( .A(A[4]), .B(B_AS[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4])
         );
  FAX1 U1_3 ( .A(A[3]), .B(B_AS[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3])
         );
  FAX1 U1_2 ( .A(A[2]), .B(B_AS[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2])
         );
  FAX1 U1_1 ( .A(A[1]), .B(B_AS[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1])
         );
  FAX1 U1_0 ( .A(A[0]), .B(B_AS[0]), .C(carry[0]), .YC(carry[1]), .YS(SUM[0])
         );
  AND2X2 U1 ( .A(n12), .B(B_AS[29]), .Y(n1) );
  AND2X2 U2 ( .A(n13), .B(B_AS[27]), .Y(n2) );
  AND2X2 U3 ( .A(n14), .B(B_AS[25]), .Y(n3) );
  AND2X2 U4 ( .A(n15), .B(B_AS[23]), .Y(n4) );
  AND2X2 U5 ( .A(n16), .B(B_AS[21]), .Y(n5) );
  AND2X2 U6 ( .A(n17), .B(B_AS[19]), .Y(n6) );
  AND2X2 U7 ( .A(n18), .B(B_AS[17]), .Y(n7) );
  AND2X2 U8 ( .A(n19), .B(B_AS[15]), .Y(n8) );
  AND2X2 U9 ( .A(n20), .B(B_AS[13]), .Y(n9) );
  AND2X2 U10 ( .A(n21), .B(B_AS[11]), .Y(n10) );
  AND2X2 U11 ( .A(n22), .B(B_AS[9]), .Y(n11) );
  AND2X2 U12 ( .A(n2), .B(B_AS[28]), .Y(n12) );
  AND2X2 U13 ( .A(n3), .B(B_AS[26]), .Y(n13) );
  AND2X2 U14 ( .A(n4), .B(B_AS[24]), .Y(n14) );
  AND2X2 U15 ( .A(n5), .B(B_AS[22]), .Y(n15) );
  AND2X2 U16 ( .A(n6), .B(B_AS[20]), .Y(n16) );
  AND2X2 U17 ( .A(n7), .B(B_AS[18]), .Y(n17) );
  AND2X2 U18 ( .A(n8), .B(B_AS[16]), .Y(n18) );
  AND2X2 U19 ( .A(n9), .B(B_AS[14]), .Y(n19) );
  AND2X2 U20 ( .A(n10), .B(B_AS[12]), .Y(n20) );
  AND2X2 U21 ( .A(n11), .B(B_AS[10]), .Y(n21) );
  AND2X2 U22 ( .A(carry[8]), .B(B_AS[8]), .Y(n22) );
  AND2X2 U23 ( .A(n1), .B(B_AS[30]), .Y(n23) );
  XOR2X1 U24 ( .A(B_AS[31]), .B(n23), .Y(SUM[31]) );
  XOR2X1 U25 ( .A(n1), .B(B_AS[30]), .Y(SUM[30]) );
  XOR2X1 U26 ( .A(n12), .B(B_AS[29]), .Y(SUM[29]) );
  XOR2X1 U27 ( .A(n2), .B(B_AS[28]), .Y(SUM[28]) );
  XOR2X1 U28 ( .A(n13), .B(B_AS[27]), .Y(SUM[27]) );
  XOR2X1 U29 ( .A(n3), .B(B_AS[26]), .Y(SUM[26]) );
  XOR2X1 U30 ( .A(n14), .B(B_AS[25]), .Y(SUM[25]) );
  XOR2X1 U31 ( .A(n4), .B(B_AS[24]), .Y(SUM[24]) );
  XOR2X1 U32 ( .A(n15), .B(B_AS[23]), .Y(SUM[23]) );
  XOR2X1 U33 ( .A(n5), .B(B_AS[22]), .Y(SUM[22]) );
  XOR2X1 U34 ( .A(n16), .B(B_AS[21]), .Y(SUM[21]) );
  XOR2X1 U35 ( .A(n6), .B(B_AS[20]), .Y(SUM[20]) );
  XOR2X1 U36 ( .A(n17), .B(B_AS[19]), .Y(SUM[19]) );
  XOR2X1 U37 ( .A(n7), .B(B_AS[18]), .Y(SUM[18]) );
  XOR2X1 U38 ( .A(n18), .B(B_AS[17]), .Y(SUM[17]) );
  XOR2X1 U39 ( .A(n8), .B(B_AS[16]), .Y(SUM[16]) );
  XOR2X1 U40 ( .A(n19), .B(B_AS[15]), .Y(SUM[15]) );
  XOR2X1 U41 ( .A(n9), .B(B_AS[14]), .Y(SUM[14]) );
  XOR2X1 U42 ( .A(n20), .B(B_AS[13]), .Y(SUM[13]) );
  XOR2X1 U43 ( .A(n10), .B(B_AS[12]), .Y(SUM[12]) );
  XOR2X1 U44 ( .A(n21), .B(B_AS[11]), .Y(SUM[11]) );
  XOR2X1 U45 ( .A(n11), .B(B_AS[10]), .Y(SUM[10]) );
  XOR2X1 U46 ( .A(n22), .B(B_AS[9]), .Y(SUM[9]) );
  XOR2X1 U47 ( .A(carry[8]), .B(B_AS[8]), .Y(SUM[8]) );
  XOR2X1 U48 ( .A(B[9]), .B(carry[0]), .Y(B_AS[9]) );
  XOR2X1 U49 ( .A(B[8]), .B(carry[0]), .Y(B_AS[8]) );
  XOR2X1 U50 ( .A(B[7]), .B(carry[0]), .Y(B_AS[7]) );
  XOR2X1 U51 ( .A(B[6]), .B(carry[0]), .Y(B_AS[6]) );
  XOR2X1 U52 ( .A(B[5]), .B(carry[0]), .Y(B_AS[5]) );
  XOR2X1 U53 ( .A(B[4]), .B(carry[0]), .Y(B_AS[4]) );
  XOR2X1 U54 ( .A(B[3]), .B(carry[0]), .Y(B_AS[3]) );
  XOR2X1 U55 ( .A(B[31]), .B(carry[0]), .Y(B_AS[31]) );
  XOR2X1 U56 ( .A(B[30]), .B(carry[0]), .Y(B_AS[30]) );
  XOR2X1 U57 ( .A(B[2]), .B(carry[0]), .Y(B_AS[2]) );
  XOR2X1 U58 ( .A(B[29]), .B(carry[0]), .Y(B_AS[29]) );
  XOR2X1 U59 ( .A(B[28]), .B(carry[0]), .Y(B_AS[28]) );
  XOR2X1 U60 ( .A(B[27]), .B(carry[0]), .Y(B_AS[27]) );
  XOR2X1 U61 ( .A(B[26]), .B(carry[0]), .Y(B_AS[26]) );
  XOR2X1 U62 ( .A(B[25]), .B(carry[0]), .Y(B_AS[25]) );
  XOR2X1 U63 ( .A(B[24]), .B(carry[0]), .Y(B_AS[24]) );
  XOR2X1 U64 ( .A(B[23]), .B(carry[0]), .Y(B_AS[23]) );
  XOR2X1 U65 ( .A(B[22]), .B(carry[0]), .Y(B_AS[22]) );
  XOR2X1 U66 ( .A(B[21]), .B(carry[0]), .Y(B_AS[21]) );
  XOR2X1 U67 ( .A(B[20]), .B(carry[0]), .Y(B_AS[20]) );
  XOR2X1 U68 ( .A(B[1]), .B(carry[0]), .Y(B_AS[1]) );
  XOR2X1 U69 ( .A(B[19]), .B(carry[0]), .Y(B_AS[19]) );
  XOR2X1 U70 ( .A(B[18]), .B(carry[0]), .Y(B_AS[18]) );
  XOR2X1 U71 ( .A(B[17]), .B(carry[0]), .Y(B_AS[17]) );
  XOR2X1 U72 ( .A(B[16]), .B(carry[0]), .Y(B_AS[16]) );
  XOR2X1 U73 ( .A(B[15]), .B(carry[0]), .Y(B_AS[15]) );
  XOR2X1 U74 ( .A(B[14]), .B(carry[0]), .Y(B_AS[14]) );
  XOR2X1 U75 ( .A(B[13]), .B(carry[0]), .Y(B_AS[13]) );
  XOR2X1 U76 ( .A(B[12]), .B(carry[0]), .Y(B_AS[12]) );
  XOR2X1 U77 ( .A(B[11]), .B(carry[0]), .Y(B_AS[11]) );
  XOR2X1 U78 ( .A(B[10]), .B(carry[0]), .Y(B_AS[10]) );
  XOR2X1 U79 ( .A(B[0]), .B(carry[0]), .Y(B_AS[0]) );
endmodule


module CannyEdge_DW01_add_48 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140;
  assign SUM[6] = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2X1 U2 ( .A(n140), .B(B[7]), .Y(SUM[7]) );
  NAND2X1 U29 ( .A(A[7]), .B(B[7]), .Y(n114) );
  XOR2X1 U30 ( .A(n28), .B(n29), .Y(SUM[9]) );
  NOR2X1 U31 ( .A(n136), .B(n30), .Y(n29) );
  XOR2X1 U32 ( .A(n32), .B(n114), .Y(SUM[8]) );
  NAND2X1 U33 ( .A(n139), .B(n33), .Y(n32) );
  XOR2X1 U34 ( .A(n35), .B(n36), .Y(SUM[29]) );
  XOR2X1 U35 ( .A(B[29]), .B(A[29]), .Y(n36) );
  OAI21X1 U36 ( .A(n37), .B(n38), .C(n39), .Y(n35) );
  XOR2X1 U37 ( .A(n40), .B(n38), .Y(SUM[28]) );
  AOI21X1 U38 ( .A(n116), .B(n41), .C(n42), .Y(n38) );
  NAND2X1 U39 ( .A(n115), .B(n39), .Y(n40) );
  NAND2X1 U40 ( .A(B[28]), .B(A[28]), .Y(n39) );
  NOR2X1 U41 ( .A(B[28]), .B(A[28]), .Y(n37) );
  XOR2X1 U42 ( .A(n41), .B(n44), .Y(SUM[27]) );
  NOR2X1 U43 ( .A(n42), .B(n43), .Y(n44) );
  NOR2X1 U44 ( .A(B[27]), .B(A[27]), .Y(n43) );
  AND2X1 U45 ( .A(B[27]), .B(A[27]), .Y(n42) );
  OAI21X1 U46 ( .A(n45), .B(n46), .C(n47), .Y(n41) );
  XOR2X1 U47 ( .A(n48), .B(n46), .Y(SUM[26]) );
  AOI21X1 U48 ( .A(n117), .B(n49), .C(n50), .Y(n46) );
  NAND2X1 U49 ( .A(n128), .B(n47), .Y(n48) );
  NAND2X1 U50 ( .A(B[26]), .B(A[26]), .Y(n47) );
  NOR2X1 U51 ( .A(B[26]), .B(A[26]), .Y(n45) );
  XOR2X1 U52 ( .A(n49), .B(n52), .Y(SUM[25]) );
  NOR2X1 U53 ( .A(n50), .B(n51), .Y(n52) );
  NOR2X1 U54 ( .A(B[25]), .B(A[25]), .Y(n51) );
  AND2X1 U55 ( .A(B[25]), .B(A[25]), .Y(n50) );
  OAI21X1 U56 ( .A(n53), .B(n54), .C(n55), .Y(n49) );
  XOR2X1 U57 ( .A(n56), .B(n54), .Y(SUM[24]) );
  AOI21X1 U58 ( .A(n119), .B(n57), .C(n58), .Y(n54) );
  NAND2X1 U59 ( .A(n118), .B(n55), .Y(n56) );
  NAND2X1 U60 ( .A(B[24]), .B(A[24]), .Y(n55) );
  NOR2X1 U61 ( .A(B[24]), .B(A[24]), .Y(n53) );
  XOR2X1 U62 ( .A(n57), .B(n60), .Y(SUM[23]) );
  NOR2X1 U63 ( .A(n58), .B(n59), .Y(n60) );
  NOR2X1 U64 ( .A(B[23]), .B(A[23]), .Y(n59) );
  AND2X1 U65 ( .A(B[23]), .B(A[23]), .Y(n58) );
  OAI21X1 U66 ( .A(n61), .B(n62), .C(n63), .Y(n57) );
  XOR2X1 U67 ( .A(n64), .B(n62), .Y(SUM[22]) );
  AOI21X1 U68 ( .A(n120), .B(n65), .C(n66), .Y(n62) );
  NAND2X1 U69 ( .A(n127), .B(n63), .Y(n64) );
  NAND2X1 U70 ( .A(B[22]), .B(A[22]), .Y(n63) );
  NOR2X1 U71 ( .A(B[22]), .B(A[22]), .Y(n61) );
  XOR2X1 U72 ( .A(n65), .B(n68), .Y(SUM[21]) );
  NOR2X1 U73 ( .A(n66), .B(n67), .Y(n68) );
  NOR2X1 U74 ( .A(B[21]), .B(A[21]), .Y(n67) );
  AND2X1 U75 ( .A(B[21]), .B(A[21]), .Y(n66) );
  OAI21X1 U76 ( .A(n69), .B(n70), .C(n71), .Y(n65) );
  XOR2X1 U77 ( .A(n72), .B(n70), .Y(SUM[20]) );
  AOI21X1 U78 ( .A(n122), .B(n73), .C(n74), .Y(n70) );
  NAND2X1 U79 ( .A(n121), .B(n71), .Y(n72) );
  NAND2X1 U80 ( .A(B[20]), .B(A[20]), .Y(n71) );
  NOR2X1 U81 ( .A(B[20]), .B(A[20]), .Y(n69) );
  XOR2X1 U82 ( .A(n73), .B(n76), .Y(SUM[19]) );
  NOR2X1 U83 ( .A(n74), .B(n75), .Y(n76) );
  NOR2X1 U84 ( .A(B[19]), .B(A[19]), .Y(n75) );
  AND2X1 U85 ( .A(B[19]), .B(A[19]), .Y(n74) );
  OAI21X1 U86 ( .A(n77), .B(n78), .C(n79), .Y(n73) );
  XOR2X1 U87 ( .A(n80), .B(n78), .Y(SUM[18]) );
  AOI21X1 U88 ( .A(n123), .B(n81), .C(n82), .Y(n78) );
  NAND2X1 U89 ( .A(n126), .B(n79), .Y(n80) );
  NAND2X1 U90 ( .A(B[18]), .B(A[18]), .Y(n79) );
  NOR2X1 U91 ( .A(B[18]), .B(A[18]), .Y(n77) );
  XOR2X1 U92 ( .A(n81), .B(n84), .Y(SUM[17]) );
  NOR2X1 U93 ( .A(n82), .B(n83), .Y(n84) );
  NOR2X1 U94 ( .A(B[17]), .B(A[17]), .Y(n83) );
  AND2X1 U95 ( .A(B[17]), .B(A[17]), .Y(n82) );
  OAI21X1 U96 ( .A(n85), .B(n86), .C(n87), .Y(n81) );
  XOR2X1 U97 ( .A(n88), .B(n86), .Y(SUM[16]) );
  AOI21X1 U98 ( .A(n125), .B(n89), .C(n90), .Y(n86) );
  NAND2X1 U99 ( .A(n124), .B(n87), .Y(n88) );
  NAND2X1 U100 ( .A(B[16]), .B(A[16]), .Y(n87) );
  NOR2X1 U101 ( .A(B[16]), .B(A[16]), .Y(n85) );
  XOR2X1 U102 ( .A(n89), .B(n92), .Y(SUM[15]) );
  NOR2X1 U103 ( .A(n90), .B(n91), .Y(n92) );
  NOR2X1 U104 ( .A(B[15]), .B(A[15]), .Y(n91) );
  AND2X1 U105 ( .A(B[15]), .B(A[15]), .Y(n90) );
  OAI21X1 U106 ( .A(n93), .B(n94), .C(n95), .Y(n89) );
  XOR2X1 U107 ( .A(n96), .B(n94), .Y(SUM[14]) );
  AOI21X1 U108 ( .A(n130), .B(n97), .C(n98), .Y(n94) );
  NAND2X1 U109 ( .A(n129), .B(n95), .Y(n96) );
  NAND2X1 U110 ( .A(B[14]), .B(A[14]), .Y(n95) );
  NOR2X1 U111 ( .A(B[14]), .B(A[14]), .Y(n93) );
  XOR2X1 U112 ( .A(n97), .B(n100), .Y(SUM[13]) );
  NOR2X1 U113 ( .A(n98), .B(n99), .Y(n100) );
  NOR2X1 U114 ( .A(B[13]), .B(A[13]), .Y(n99) );
  AND2X1 U115 ( .A(B[13]), .B(A[13]), .Y(n98) );
  OAI21X1 U116 ( .A(n101), .B(n132), .C(n102), .Y(n97) );
  XOR2X1 U117 ( .A(n103), .B(n132), .Y(SUM[12]) );
  OAI21X1 U118 ( .A(n105), .B(n106), .C(n107), .Y(n104) );
  AOI21X1 U119 ( .A(n108), .B(n135), .C(n134), .Y(n106) );
  NAND2X1 U120 ( .A(n131), .B(n102), .Y(n103) );
  NAND2X1 U121 ( .A(B[12]), .B(A[12]), .Y(n102) );
  NOR2X1 U122 ( .A(B[12]), .B(A[12]), .Y(n101) );
  XOR2X1 U123 ( .A(n110), .B(n111), .Y(SUM[11]) );
  NOR2X1 U124 ( .A(n133), .B(n105), .Y(n111) );
  NOR2X1 U125 ( .A(B[11]), .B(A[11]), .Y(n105) );
  NAND2X1 U126 ( .A(B[11]), .B(A[11]), .Y(n107) );
  OAI21X1 U127 ( .A(n112), .B(n137), .C(n109), .Y(n110) );
  XOR2X1 U128 ( .A(n113), .B(n137), .Y(SUM[10]) );
  OAI21X1 U129 ( .A(n138), .B(n30), .C(n31), .Y(n108) );
  NAND2X1 U130 ( .A(B[9]), .B(A[9]), .Y(n31) );
  NOR2X1 U131 ( .A(B[9]), .B(A[9]), .Y(n30) );
  OAI21X1 U132 ( .A(n34), .B(n114), .C(n33), .Y(n28) );
  NAND2X1 U133 ( .A(B[8]), .B(A[8]), .Y(n33) );
  NOR2X1 U134 ( .A(B[8]), .B(A[8]), .Y(n34) );
  NAND2X1 U135 ( .A(n135), .B(n109), .Y(n113) );
  NAND2X1 U136 ( .A(B[10]), .B(A[10]), .Y(n109) );
  NOR2X1 U137 ( .A(B[10]), .B(A[10]), .Y(n112) );
  INVX2 U3 ( .A(n37), .Y(n115) );
  INVX2 U4 ( .A(n43), .Y(n116) );
  INVX2 U5 ( .A(n51), .Y(n117) );
  INVX2 U6 ( .A(n53), .Y(n118) );
  INVX2 U7 ( .A(n59), .Y(n119) );
  INVX2 U8 ( .A(n67), .Y(n120) );
  INVX2 U9 ( .A(n69), .Y(n121) );
  INVX2 U10 ( .A(n75), .Y(n122) );
  INVX2 U11 ( .A(n83), .Y(n123) );
  INVX2 U12 ( .A(n85), .Y(n124) );
  INVX2 U13 ( .A(n91), .Y(n125) );
  INVX2 U14 ( .A(n77), .Y(n126) );
  INVX2 U15 ( .A(n61), .Y(n127) );
  INVX2 U16 ( .A(n45), .Y(n128) );
  INVX2 U17 ( .A(n93), .Y(n129) );
  INVX2 U18 ( .A(n99), .Y(n130) );
  INVX2 U19 ( .A(n101), .Y(n131) );
  INVX2 U20 ( .A(n104), .Y(n132) );
  INVX2 U21 ( .A(n107), .Y(n133) );
  INVX2 U22 ( .A(n109), .Y(n134) );
  INVX2 U23 ( .A(n112), .Y(n135) );
  INVX2 U24 ( .A(n31), .Y(n136) );
  INVX2 U25 ( .A(n108), .Y(n137) );
  INVX2 U26 ( .A(n28), .Y(n138) );
  INVX2 U27 ( .A(n34), .Y(n139) );
  INVX2 U28 ( .A(A[7]), .Y(n140) );
endmodule


module CannyEdge_DW02_mult_24 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [31:0] B;
  output [39:0] PRODUCT;
  input TC;
  wire   \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \CARRYB[7][0] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[7][1] ,
         \SUMB[7][0] , \SUMB[6][1] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] ,
         \SUMB[3][1] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] ,
         \SUMB[2][1] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[36] , \A1[35] , \A1[34] , \A1[33] ,
         \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] ,
         \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[4] ,
         \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n130, n131, n132, n133, n134, n135, n136,
         n137, n145, n143, n142, n141, n140, n139, n138, n129, n12, n114,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][30] , \SUMB[7][2] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][30] , \SUMB[6][2] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][30] , \SUMB[5][29] ,
         \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] , \SUMB[5][25] ,
         \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] ,
         \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] ,
         \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] ,
         \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] , \SUMB[4][9] ,
         \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][30] , \SUMB[3][29] , \SUMB[3][28] ,
         \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] ,
         \SUMB[3][23] , \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] ,
         \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] , \SUMB[3][16] ,
         \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] ,
         \SUMB[3][11] , \SUMB[3][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][30] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[1][7] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][30] ,
         \CARRYB[7][2] , \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] ,
         \CARRYB[7][26] , \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] ,
         \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][1] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][30] , \CARRYB[6][2] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][30] , \CARRYB[5][29] ,
         \CARRYB[5][28] , \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] ,
         \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][30] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][30] , \CARRYB[2][29] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n144, n146, n147,
         n148, n149, n150, n151, n152, n153, n154;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  FAX1 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .C(\SUMB[6][1] ), .YC(
        \CARRYB[7][0] ), .YS(\SUMB[7][0] ) );
  FAX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .C(\SUMB[5][1] ), .YC(
        \CARRYB[6][0] ), .YS(\A1[4] ) );
  FAX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .C(\SUMB[5][2] ), .YC(
        \CARRYB[6][1] ), .YS(\SUMB[6][1] ) );
  FAX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .C(\SUMB[4][1] ), .YC(
        \CARRYB[5][0] ), .YS(\A1[3] ) );
  FAX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .C(\SUMB[4][2] ), .YC(
        \CARRYB[5][1] ), .YS(\SUMB[5][1] ) );
  FAX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .C(\SUMB[4][3] ), .YC(
        \CARRYB[5][2] ), .YS(\SUMB[5][2] ) );
  FAX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .C(\SUMB[3][1] ), .YC(
        \CARRYB[4][0] ), .YS(\A1[2] ) );
  FAX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .C(\SUMB[3][2] ), .YC(
        \CARRYB[4][1] ), .YS(\SUMB[4][1] ) );
  FAX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .C(\SUMB[3][3] ), .YC(
        \CARRYB[4][2] ), .YS(\SUMB[4][2] ) );
  FAX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .C(\SUMB[3][4] ), .YC(
        \CARRYB[4][3] ), .YS(\SUMB[4][3] ) );
  FAX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .C(\SUMB[2][1] ), .YC(
        \CARRYB[3][0] ), .YS(\A1[1] ) );
  FAX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .C(\SUMB[2][2] ), .YC(
        \CARRYB[3][1] ), .YS(\SUMB[3][1] ) );
  FAX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .C(\SUMB[2][3] ), .YC(
        \CARRYB[3][2] ), .YS(\SUMB[3][2] ) );
  FAX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .C(\SUMB[2][4] ), .YC(
        \CARRYB[3][3] ), .YS(\SUMB[3][3] ) );
  FAX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .C(\SUMB[2][5] ), .YC(
        \CARRYB[3][4] ), .YS(\SUMB[3][4] ) );
  FAX1 S1_2_0 ( .A(\ab[2][0] ), .B(n19), .C(\SUMB[1][1] ), .YC(\CARRYB[2][0] ), 
        .YS(\A1[0] ) );
  FAX1 S2_2_1 ( .A(\ab[2][1] ), .B(n18), .C(\SUMB[1][2] ), .YC(\CARRYB[2][1] ), 
        .YS(\SUMB[2][1] ) );
  FAX1 S2_2_2 ( .A(\ab[2][2] ), .B(n17), .C(\SUMB[1][3] ), .YC(\CARRYB[2][2] ), 
        .YS(\SUMB[2][2] ) );
  FAX1 S2_2_3 ( .A(\ab[2][3] ), .B(n16), .C(\SUMB[1][4] ), .YC(\CARRYB[2][3] ), 
        .YS(\SUMB[2][3] ) );
  FAX1 S2_2_4 ( .A(\ab[2][4] ), .B(n15), .C(\SUMB[1][5] ), .YC(\CARRYB[2][4] ), 
        .YS(\SUMB[2][4] ) );
  FAX1 S2_2_5 ( .A(\ab[2][5] ), .B(n14), .C(\SUMB[1][6] ), .YC(\CARRYB[2][5] ), 
        .YS(\SUMB[2][5] ) );
  OR2X2 U5 ( .A(n116), .B(n109), .Y(n115) );
  OR2X2 U6 ( .A(n118), .B(n109), .Y(n117) );
  OR2X2 U7 ( .A(n120), .B(n109), .Y(n119) );
  OR2X2 U8 ( .A(n122), .B(n109), .Y(n121) );
  OR2X2 U9 ( .A(n124), .B(n109), .Y(n123) );
  OR2X2 U10 ( .A(n126), .B(n109), .Y(n125) );
  OR2X2 U11 ( .A(n128), .B(n109), .Y(n127) );
  AND2X1 U64 ( .A(\CARRYB[7][0] ), .B(\SUMB[7][1] ), .Y(n20) );
  NOR2X1 U65 ( .A(n148), .B(n115), .Y(n19) );
  NOR2X1 U66 ( .A(n149), .B(n117), .Y(n18) );
  NOR2X1 U67 ( .A(n150), .B(n119), .Y(n17) );
  NOR2X1 U68 ( .A(n151), .B(n121), .Y(n16) );
  NOR2X1 U69 ( .A(n152), .B(n123), .Y(n15) );
  NOR2X1 U70 ( .A(n153), .B(n125), .Y(n14) );
  NOR2X1 U71 ( .A(n154), .B(n127), .Y(n13) );
  NOR2X1 U75 ( .A(n146), .B(n154), .Y(\ab[7][7] ) );
  NOR2X1 U76 ( .A(n146), .B(n153), .Y(\ab[7][6] ) );
  NOR2X1 U77 ( .A(n146), .B(n152), .Y(\ab[7][5] ) );
  NOR2X1 U78 ( .A(n146), .B(n151), .Y(\ab[7][4] ) );
  NOR2X1 U79 ( .A(n146), .B(n150), .Y(\ab[7][3] ) );
  NOR2X1 U80 ( .A(n146), .B(n149), .Y(\ab[7][2] ) );
  NOR2X1 U81 ( .A(n146), .B(n148), .Y(\ab[7][1] ) );
  NOR2X1 U82 ( .A(n146), .B(n147), .Y(\ab[7][0] ) );
  NOR2X1 U83 ( .A(n144), .B(n154), .Y(\ab[6][7] ) );
  NOR2X1 U84 ( .A(n144), .B(n153), .Y(\ab[6][6] ) );
  NOR2X1 U85 ( .A(n144), .B(n152), .Y(\ab[6][5] ) );
  NOR2X1 U86 ( .A(n144), .B(n151), .Y(\ab[6][4] ) );
  NOR2X1 U87 ( .A(n144), .B(n150), .Y(\ab[6][3] ) );
  NOR2X1 U88 ( .A(n144), .B(n149), .Y(\ab[6][2] ) );
  NOR2X1 U89 ( .A(n144), .B(n148), .Y(\ab[6][1] ) );
  NOR2X1 U90 ( .A(n144), .B(n147), .Y(\ab[6][0] ) );
  NOR2X1 U91 ( .A(n113), .B(n154), .Y(\ab[5][7] ) );
  NOR2X1 U92 ( .A(n113), .B(n153), .Y(\ab[5][6] ) );
  NOR2X1 U93 ( .A(n113), .B(n152), .Y(\ab[5][5] ) );
  NOR2X1 U94 ( .A(n113), .B(n151), .Y(\ab[5][4] ) );
  NOR2X1 U95 ( .A(n113), .B(n150), .Y(\ab[5][3] ) );
  NOR2X1 U96 ( .A(n113), .B(n149), .Y(\ab[5][2] ) );
  NOR2X1 U97 ( .A(n113), .B(n148), .Y(\ab[5][1] ) );
  NOR2X1 U98 ( .A(n113), .B(n147), .Y(\ab[5][0] ) );
  NOR2X1 U99 ( .A(n112), .B(n154), .Y(\ab[4][7] ) );
  NOR2X1 U100 ( .A(n112), .B(n153), .Y(\ab[4][6] ) );
  NOR2X1 U101 ( .A(n112), .B(n152), .Y(\ab[4][5] ) );
  NOR2X1 U102 ( .A(n112), .B(n151), .Y(\ab[4][4] ) );
  NOR2X1 U103 ( .A(n112), .B(n150), .Y(\ab[4][3] ) );
  NOR2X1 U104 ( .A(n112), .B(n149), .Y(\ab[4][2] ) );
  NOR2X1 U105 ( .A(n112), .B(n148), .Y(\ab[4][1] ) );
  NOR2X1 U106 ( .A(n112), .B(n147), .Y(\ab[4][0] ) );
  NOR2X1 U107 ( .A(n111), .B(n154), .Y(\ab[3][7] ) );
  NOR2X1 U108 ( .A(n111), .B(n153), .Y(\ab[3][6] ) );
  NOR2X1 U109 ( .A(n111), .B(n152), .Y(\ab[3][5] ) );
  NOR2X1 U110 ( .A(n111), .B(n151), .Y(\ab[3][4] ) );
  NOR2X1 U111 ( .A(n111), .B(n150), .Y(\ab[3][3] ) );
  NOR2X1 U112 ( .A(n111), .B(n149), .Y(\ab[3][2] ) );
  NOR2X1 U113 ( .A(n111), .B(n148), .Y(\ab[3][1] ) );
  NOR2X1 U114 ( .A(n111), .B(n147), .Y(\ab[3][0] ) );
  NOR2X1 U115 ( .A(n110), .B(n154), .Y(\ab[2][7] ) );
  NOR2X1 U116 ( .A(n110), .B(n153), .Y(\ab[2][6] ) );
  NOR2X1 U117 ( .A(n110), .B(n152), .Y(\ab[2][5] ) );
  NOR2X1 U118 ( .A(n110), .B(n151), .Y(\ab[2][4] ) );
  NOR2X1 U119 ( .A(n110), .B(n150), .Y(\ab[2][3] ) );
  NOR2X1 U120 ( .A(n110), .B(n149), .Y(\ab[2][2] ) );
  NOR2X1 U121 ( .A(n110), .B(n148), .Y(\ab[2][1] ) );
  NOR2X1 U122 ( .A(n110), .B(n147), .Y(\ab[2][0] ) );
  NAND2X1 U124 ( .A(B[7]), .B(A[1]), .Y(n130) );
  XOR2X1 U125 ( .A(n128), .B(n131), .Y(\SUMB[1][6] ) );
  NAND2X1 U126 ( .A(B[7]), .B(A[0]), .Y(n131) );
  NAND2X1 U127 ( .A(B[6]), .B(A[1]), .Y(n128) );
  XOR2X1 U128 ( .A(n126), .B(n132), .Y(\SUMB[1][5] ) );
  NAND2X1 U129 ( .A(B[6]), .B(A[0]), .Y(n132) );
  NAND2X1 U130 ( .A(B[5]), .B(A[1]), .Y(n126) );
  XOR2X1 U131 ( .A(n124), .B(n133), .Y(\SUMB[1][4] ) );
  NAND2X1 U132 ( .A(B[5]), .B(A[0]), .Y(n133) );
  NAND2X1 U133 ( .A(B[4]), .B(A[1]), .Y(n124) );
  XOR2X1 U134 ( .A(n122), .B(n134), .Y(\SUMB[1][3] ) );
  NAND2X1 U135 ( .A(B[4]), .B(A[0]), .Y(n134) );
  NAND2X1 U136 ( .A(B[3]), .B(A[1]), .Y(n122) );
  XOR2X1 U137 ( .A(n120), .B(n135), .Y(\SUMB[1][2] ) );
  NAND2X1 U138 ( .A(B[3]), .B(A[0]), .Y(n135) );
  NAND2X1 U139 ( .A(B[2]), .B(A[1]), .Y(n120) );
  XOR2X1 U140 ( .A(n118), .B(n136), .Y(\SUMB[1][1] ) );
  NAND2X1 U141 ( .A(B[2]), .B(A[0]), .Y(n136) );
  NAND2X1 U142 ( .A(B[1]), .B(A[1]), .Y(n118) );
  XOR2X1 U146 ( .A(n116), .B(n137), .Y(PRODUCT[1]) );
  NAND2X1 U147 ( .A(B[1]), .B(A[0]), .Y(n137) );
  NAND2X1 U148 ( .A(B[0]), .B(A[1]), .Y(n116) );
  NOR2X1 U149 ( .A(n109), .B(n147), .Y(PRODUCT[0]) );
  XOR2X1 U153 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Y(\A1[6] ) );
  CannyEdge_DW01_add_48 FS_1 ( .A({1'b0, \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \SUMB[7][0] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({n3, 
        n4, n5, n6, n7, n8, n9, n10, n21, n29, n22, n30, n23, n31, n24, n32, 
        n25, n33, n26, n34, n27, n35, n28, n37, n36, n38, n39, n42, n40, n41, 
        n20, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, PRODUCT[31:2]}) );
  XOR2X1 U154 ( .A(\CARRYB[7][30] ), .B(n106), .Y(\A1[36] ) );
  AND2X1 U54 ( .A(n106), .B(\CARRYB[7][30] ), .Y(n3) );
  XOR2X1 U152 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Y(\A1[7] ) );
  AND2X1 U41 ( .A(\CARRYB[7][1] ), .B(\SUMB[7][2] ), .Y(n41) );
  FAX1 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .C(\SUMB[6][2] ), .YC(
        \CARRYB[7][1] ), .YS(\SUMB[7][1] ) );
  XOR2X1 U151 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Y(\A1[8] ) );
  AND2X1 U42 ( .A(\CARRYB[7][2] ), .B(\SUMB[7][3] ), .Y(n40) );
  FAX1 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .C(\SUMB[6][3] ), .YC(
        \CARRYB[7][2] ), .YS(\SUMB[7][2] ) );
  FAX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .C(\SUMB[5][3] ), .YC(
        \CARRYB[6][2] ), .YS(\SUMB[6][2] ) );
  XOR2X1 U150 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Y(\A1[9] ) );
  AND2X1 U40 ( .A(\CARRYB[7][3] ), .B(\SUMB[7][4] ), .Y(n42) );
  FAX1 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .C(\SUMB[6][4] ), .YC(
        \CARRYB[7][3] ), .YS(\SUMB[7][3] ) );
  FAX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .C(\SUMB[5][4] ), .YC(
        \CARRYB[6][3] ), .YS(\SUMB[6][3] ) );
  FAX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .C(\SUMB[4][4] ), .YC(
        \CARRYB[5][3] ), .YS(\SUMB[5][3] ) );
  XOR2X1 U181 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Y(\A1[10] ) );
  AND2X1 U44 ( .A(\CARRYB[7][4] ), .B(\SUMB[7][5] ), .Y(n39) );
  FAX1 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .C(\SUMB[6][5] ), .YC(
        \CARRYB[7][4] ), .YS(\SUMB[7][4] ) );
  FAX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .C(\SUMB[5][5] ), .YC(
        \CARRYB[6][4] ), .YS(\SUMB[6][4] ) );
  FAX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .C(\SUMB[4][5] ), .YC(
        \CARRYB[5][4] ), .YS(\SUMB[5][4] ) );
  FAX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .C(\SUMB[3][5] ), .YC(
        \CARRYB[4][4] ), .YS(\SUMB[4][4] ) );
  XOR2X1 U180 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Y(\A1[11] ) );
  AND2X1 U45 ( .A(\CARRYB[7][5] ), .B(\SUMB[7][6] ), .Y(n38) );
  FAX1 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .C(\SUMB[6][6] ), .YC(
        \CARRYB[7][5] ), .YS(\SUMB[7][5] ) );
  FAX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .C(\SUMB[5][6] ), .YC(
        \CARRYB[6][5] ), .YS(\SUMB[6][5] ) );
  FAX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .C(\SUMB[4][6] ), .YC(
        \CARRYB[5][5] ), .YS(\SUMB[5][5] ) );
  FAX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .C(\SUMB[3][6] ), .YC(
        \CARRYB[4][5] ), .YS(\SUMB[4][5] ) );
  FAX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .C(\SUMB[2][6] ), .YC(
        \CARRYB[3][5] ), .YS(\SUMB[3][5] ) );
  XOR2X1 U179 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Y(\A1[12] ) );
  AND2X1 U47 ( .A(\CARRYB[7][6] ), .B(\SUMB[7][7] ), .Y(n36) );
  FAX1 S4_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .C(\SUMB[6][7] ), .YC(
        \CARRYB[7][6] ), .YS(\SUMB[7][6] ) );
  FAX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .C(\SUMB[5][7] ), .YC(
        \CARRYB[6][6] ), .YS(\SUMB[6][6] ) );
  FAX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .C(\SUMB[4][7] ), .YC(
        \CARRYB[5][6] ), .YS(\SUMB[5][6] ) );
  FAX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .C(\SUMB[3][7] ), .YC(
        \CARRYB[4][6] ), .YS(\SUMB[4][6] ) );
  FAX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .C(\SUMB[2][7] ), .YC(
        \CARRYB[3][6] ), .YS(\SUMB[3][6] ) );
  FAX1 S2_2_6 ( .A(\ab[2][6] ), .B(n13), .C(\SUMB[1][7] ), .YC(\CARRYB[2][6] ), 
        .YS(\SUMB[2][6] ) );
  XNOR2X1 U123 ( .A(n114), .B(n130), .Y(\SUMB[1][7] ) );
  XOR2X1 U175 ( .A(\SUMB[7][11] ), .B(\CARRYB[7][10] ), .Y(\A1[16] ) );
  AND2X1 U57 ( .A(\CARRYB[7][10] ), .B(\SUMB[7][11] ), .Y(n27) );
  XOR2X1 U174 ( .A(\SUMB[7][12] ), .B(\CARRYB[7][11] ), .Y(\A1[17] ) );
  AND2X1 U49 ( .A(\CARRYB[7][11] ), .B(\SUMB[7][12] ), .Y(n34) );
  FAX1 S4_11 ( .A(n106), .B(\CARRYB[6][11] ), .C(\SUMB[6][12] ), .YC(
        \CARRYB[7][11] ), .YS(\SUMB[7][11] ) );
  XOR2X1 U171 ( .A(\SUMB[7][15] ), .B(\CARRYB[7][14] ), .Y(\A1[20] ) );
  AND2X1 U59 ( .A(\CARRYB[7][14] ), .B(\SUMB[7][15] ), .Y(n25) );
  XOR2X1 U170 ( .A(\SUMB[7][16] ), .B(\CARRYB[7][15] ), .Y(\A1[21] ) );
  AND2X1 U51 ( .A(\CARRYB[7][15] ), .B(\SUMB[7][16] ), .Y(n32) );
  FAX1 S4_15 ( .A(n106), .B(\CARRYB[6][15] ), .C(\SUMB[6][16] ), .YC(
        \CARRYB[7][15] ), .YS(\SUMB[7][15] ) );
  XOR2X1 U167 ( .A(\SUMB[7][19] ), .B(\CARRYB[7][18] ), .Y(\A1[24] ) );
  AND2X1 U61 ( .A(\CARRYB[7][18] ), .B(\SUMB[7][19] ), .Y(n23) );
  XOR2X1 U166 ( .A(\SUMB[7][20] ), .B(\CARRYB[7][19] ), .Y(\A1[25] ) );
  AND2X1 U53 ( .A(\CARRYB[7][19] ), .B(\SUMB[7][20] ), .Y(n30) );
  FAX1 S4_19 ( .A(n106), .B(\CARRYB[6][19] ), .C(\SUMB[6][20] ), .YC(
        \CARRYB[7][19] ), .YS(\SUMB[7][19] ) );
  XOR2X1 U163 ( .A(\SUMB[7][23] ), .B(\CARRYB[7][22] ), .Y(\A1[28] ) );
  AND2X1 U63 ( .A(\CARRYB[7][22] ), .B(\SUMB[7][23] ), .Y(n21) );
  XOR2X1 U162 ( .A(\SUMB[7][24] ), .B(\CARRYB[7][23] ), .Y(\A1[29] ) );
  AND2X1 U74 ( .A(\CARRYB[7][23] ), .B(\SUMB[7][24] ), .Y(n10) );
  FAX1 S4_23 ( .A(n106), .B(\CARRYB[6][23] ), .C(\SUMB[6][24] ), .YC(
        \CARRYB[7][23] ), .YS(\SUMB[7][23] ) );
  XOR2X1 U159 ( .A(\SUMB[7][27] ), .B(\CARRYB[7][26] ), .Y(\A1[32] ) );
  AND2X1 U37 ( .A(\CARRYB[7][26] ), .B(\SUMB[7][27] ), .Y(n7) );
  XOR2X1 U158 ( .A(\SUMB[7][28] ), .B(\CARRYB[7][27] ), .Y(\A1[33] ) );
  AND2X1 U38 ( .A(\CARRYB[7][27] ), .B(\SUMB[7][28] ), .Y(n6) );
  FAX1 S4_27 ( .A(n106), .B(\CARRYB[6][27] ), .C(\SUMB[6][28] ), .YC(
        \CARRYB[7][27] ), .YS(\SUMB[7][27] ) );
  XOR2X1 U178 ( .A(\SUMB[7][8] ), .B(\CARRYB[7][7] ), .Y(\A1[13] ) );
  AND2X1 U46 ( .A(\CARRYB[7][7] ), .B(\SUMB[7][8] ), .Y(n37) );
  FAX1 S4_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .C(\SUMB[6][8] ), .YC(
        \CARRYB[7][7] ), .YS(\SUMB[7][7] ) );
  FAX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .C(\SUMB[5][8] ), .YC(
        \CARRYB[6][7] ), .YS(\SUMB[6][7] ) );
  FAX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .C(\SUMB[4][8] ), .YC(
        \CARRYB[5][7] ), .YS(\SUMB[5][7] ) );
  FAX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .C(\SUMB[3][8] ), .YC(
        \CARRYB[4][7] ), .YS(\SUMB[4][7] ) );
  FAX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .C(\SUMB[2][8] ), .YC(
        \CARRYB[3][7] ), .YS(\SUMB[3][7] ) );
  FAX1 S2_2_7 ( .A(\ab[2][7] ), .B(n12), .C(n101), .YC(\CARRYB[2][7] ), .YS(
        \SUMB[2][7] ) );
  NOR2X1 U72 ( .A(n154), .B(n129), .Y(n12) );
  NAND2X1 U73 ( .A(n114), .B(A[1]), .Y(n129) );
  XOR2X1 U177 ( .A(\SUMB[7][9] ), .B(\CARRYB[7][8] ), .Y(\A1[14] ) );
  AND2X1 U56 ( .A(\CARRYB[7][8] ), .B(\SUMB[7][9] ), .Y(n28) );
  FAX1 S4_8 ( .A(n106), .B(\CARRYB[6][8] ), .C(\SUMB[6][9] ), .YC(
        \CARRYB[7][8] ), .YS(\SUMB[7][8] ) );
  FAX1 S2_6_8 ( .A(n97), .B(\CARRYB[5][8] ), .C(\SUMB[5][9] ), .YC(
        \CARRYB[6][8] ), .YS(\SUMB[6][8] ) );
  FAX1 S2_5_8 ( .A(n98), .B(\CARRYB[4][8] ), .C(\SUMB[4][9] ), .YC(
        \CARRYB[5][8] ), .YS(\SUMB[5][8] ) );
  FAX1 S2_4_8 ( .A(n99), .B(\CARRYB[3][8] ), .C(\SUMB[3][9] ), .YC(
        \CARRYB[4][8] ), .YS(\SUMB[4][8] ) );
  FAX1 S2_3_8 ( .A(n102), .B(\CARRYB[2][8] ), .C(\SUMB[2][9] ), .YC(
        \CARRYB[3][8] ), .YS(\SUMB[3][8] ) );
  FAX1 S2_2_8 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][8] ), .YS(
        \SUMB[2][8] ) );
  XOR2X1 U157 ( .A(\SUMB[7][29] ), .B(\CARRYB[7][28] ), .Y(\A1[34] ) );
  AND2X1 U39 ( .A(\CARRYB[7][28] ), .B(\SUMB[7][29] ), .Y(n5) );
  FAX1 S4_28 ( .A(n106), .B(\CARRYB[6][28] ), .C(\SUMB[6][29] ), .YC(
        \CARRYB[7][28] ), .YS(\SUMB[7][28] ) );
  FAX1 S2_6_28 ( .A(n97), .B(\CARRYB[5][28] ), .C(\SUMB[5][29] ), .YC(
        \CARRYB[6][28] ), .YS(\SUMB[6][28] ) );
  XOR2X1 U161 ( .A(\SUMB[7][25] ), .B(\CARRYB[7][24] ), .Y(\A1[30] ) );
  AND2X1 U35 ( .A(\CARRYB[7][24] ), .B(\SUMB[7][25] ), .Y(n9) );
  FAX1 S4_24 ( .A(n106), .B(\CARRYB[6][24] ), .C(\SUMB[6][25] ), .YC(
        \CARRYB[7][24] ), .YS(\SUMB[7][24] ) );
  FAX1 S2_6_24 ( .A(n97), .B(\CARRYB[5][24] ), .C(\SUMB[5][25] ), .YC(
        \CARRYB[6][24] ), .YS(\SUMB[6][24] ) );
  XOR2X1 U165 ( .A(\SUMB[7][21] ), .B(\CARRYB[7][20] ), .Y(\A1[26] ) );
  AND2X1 U62 ( .A(\CARRYB[7][20] ), .B(\SUMB[7][21] ), .Y(n22) );
  FAX1 S4_20 ( .A(n106), .B(\CARRYB[6][20] ), .C(\SUMB[6][21] ), .YC(
        \CARRYB[7][20] ), .YS(\SUMB[7][20] ) );
  FAX1 S2_6_20 ( .A(n97), .B(\CARRYB[5][20] ), .C(\SUMB[5][21] ), .YC(
        \CARRYB[6][20] ), .YS(\SUMB[6][20] ) );
  XOR2X1 U169 ( .A(\SUMB[7][17] ), .B(\CARRYB[7][16] ), .Y(\A1[22] ) );
  AND2X1 U60 ( .A(\CARRYB[7][16] ), .B(\SUMB[7][17] ), .Y(n24) );
  FAX1 S4_16 ( .A(n106), .B(\CARRYB[6][16] ), .C(\SUMB[6][17] ), .YC(
        \CARRYB[7][16] ), .YS(\SUMB[7][16] ) );
  FAX1 S2_6_16 ( .A(n97), .B(\CARRYB[5][16] ), .C(\SUMB[5][17] ), .YC(
        \CARRYB[6][16] ), .YS(\SUMB[6][16] ) );
  XOR2X1 U173 ( .A(\SUMB[7][13] ), .B(\CARRYB[7][12] ), .Y(\A1[18] ) );
  AND2X1 U58 ( .A(\CARRYB[7][12] ), .B(\SUMB[7][13] ), .Y(n26) );
  FAX1 S4_12 ( .A(n106), .B(\CARRYB[6][12] ), .C(\SUMB[6][13] ), .YC(
        \CARRYB[7][12] ), .YS(\SUMB[7][12] ) );
  FAX1 S2_6_12 ( .A(n97), .B(\CARRYB[5][12] ), .C(\SUMB[5][13] ), .YC(
        \CARRYB[6][12] ), .YS(\SUMB[6][12] ) );
  XOR2X1 U176 ( .A(\SUMB[7][10] ), .B(\CARRYB[7][9] ), .Y(\A1[15] ) );
  AND2X1 U48 ( .A(\CARRYB[7][9] ), .B(\SUMB[7][10] ), .Y(n35) );
  FAX1 S4_10 ( .A(n106), .B(\CARRYB[6][10] ), .C(\SUMB[6][11] ), .YC(
        \CARRYB[7][10] ), .YS(\SUMB[7][10] ) );
  FAX1 S2_6_11 ( .A(n97), .B(\CARRYB[5][11] ), .C(\SUMB[5][12] ), .YC(
        \CARRYB[6][11] ), .YS(\SUMB[6][11] ) );
  FAX1 S2_5_12 ( .A(n98), .B(\CARRYB[4][12] ), .C(\SUMB[4][13] ), .YC(
        \CARRYB[5][12] ), .YS(\SUMB[5][12] ) );
  FAX1 S4_9 ( .A(n106), .B(\CARRYB[6][9] ), .C(\SUMB[6][10] ), .YC(
        \CARRYB[7][9] ), .YS(\SUMB[7][9] ) );
  FAX1 S2_6_10 ( .A(n97), .B(\CARRYB[5][10] ), .C(\SUMB[5][11] ), .YC(
        \CARRYB[6][10] ), .YS(\SUMB[6][10] ) );
  FAX1 S2_5_11 ( .A(n98), .B(\CARRYB[4][11] ), .C(\SUMB[4][12] ), .YC(
        \CARRYB[5][11] ), .YS(\SUMB[5][11] ) );
  FAX1 S2_4_12 ( .A(n99), .B(\CARRYB[3][12] ), .C(\SUMB[3][13] ), .YC(
        \CARRYB[4][12] ), .YS(\SUMB[4][12] ) );
  FAX1 S2_6_9 ( .A(n97), .B(\CARRYB[5][9] ), .C(\SUMB[5][10] ), .YC(
        \CARRYB[6][9] ), .YS(\SUMB[6][9] ) );
  FAX1 S2_5_10 ( .A(n98), .B(\CARRYB[4][10] ), .C(\SUMB[4][11] ), .YC(
        \CARRYB[5][10] ), .YS(\SUMB[5][10] ) );
  FAX1 S2_4_11 ( .A(n99), .B(\CARRYB[3][11] ), .C(\SUMB[3][12] ), .YC(
        \CARRYB[4][11] ), .YS(\SUMB[4][11] ) );
  FAX1 S2_3_12 ( .A(n102), .B(\CARRYB[2][12] ), .C(\SUMB[2][13] ), .YC(
        \CARRYB[3][12] ), .YS(\SUMB[3][12] ) );
  FAX1 S2_5_9 ( .A(n98), .B(\CARRYB[4][9] ), .C(\SUMB[4][10] ), .YC(
        \CARRYB[5][9] ), .YS(\SUMB[5][9] ) );
  FAX1 S2_4_10 ( .A(n99), .B(\CARRYB[3][10] ), .C(\SUMB[3][11] ), .YC(
        \CARRYB[4][10] ), .YS(\SUMB[4][10] ) );
  FAX1 S2_3_11 ( .A(n102), .B(\CARRYB[2][11] ), .C(\SUMB[2][12] ), .YC(
        \CARRYB[3][11] ), .YS(\SUMB[3][11] ) );
  FAX1 S2_2_12 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][12] ), .YS(
        \SUMB[2][12] ) );
  FAX1 S2_4_9 ( .A(n99), .B(\CARRYB[3][9] ), .C(\SUMB[3][10] ), .YC(
        \CARRYB[4][9] ), .YS(\SUMB[4][9] ) );
  FAX1 S2_3_10 ( .A(n102), .B(\CARRYB[2][10] ), .C(\SUMB[2][11] ), .YC(
        \CARRYB[3][10] ), .YS(\SUMB[3][10] ) );
  FAX1 S2_2_11 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][11] ), .YS(
        \SUMB[2][11] ) );
  FAX1 S2_3_9 ( .A(n102), .B(\CARRYB[2][9] ), .C(\SUMB[2][10] ), .YC(
        \CARRYB[3][9] ), .YS(\SUMB[3][9] ) );
  FAX1 S2_2_10 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][10] ), .YS(
        \SUMB[2][10] ) );
  FAX1 S2_2_9 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][9] ), .YS(
        \SUMB[2][9] ) );
  XOR2X1 U172 ( .A(\SUMB[7][14] ), .B(\CARRYB[7][13] ), .Y(\A1[19] ) );
  AND2X1 U50 ( .A(\CARRYB[7][13] ), .B(\SUMB[7][14] ), .Y(n33) );
  FAX1 S4_14 ( .A(n106), .B(\CARRYB[6][14] ), .C(\SUMB[6][15] ), .YC(
        \CARRYB[7][14] ), .YS(\SUMB[7][14] ) );
  FAX1 S2_6_15 ( .A(n97), .B(\CARRYB[5][15] ), .C(\SUMB[5][16] ), .YC(
        \CARRYB[6][15] ), .YS(\SUMB[6][15] ) );
  FAX1 S2_5_16 ( .A(n98), .B(\CARRYB[4][16] ), .C(\SUMB[4][17] ), .YC(
        \CARRYB[5][16] ), .YS(\SUMB[5][16] ) );
  FAX1 S4_13 ( .A(n106), .B(\CARRYB[6][13] ), .C(\SUMB[6][14] ), .YC(
        \CARRYB[7][13] ), .YS(\SUMB[7][13] ) );
  FAX1 S2_6_14 ( .A(n97), .B(\CARRYB[5][14] ), .C(\SUMB[5][15] ), .YC(
        \CARRYB[6][14] ), .YS(\SUMB[6][14] ) );
  FAX1 S2_5_15 ( .A(n98), .B(\CARRYB[4][15] ), .C(\SUMB[4][16] ), .YC(
        \CARRYB[5][15] ), .YS(\SUMB[5][15] ) );
  FAX1 S2_4_16 ( .A(n99), .B(\CARRYB[3][16] ), .C(\SUMB[3][17] ), .YC(
        \CARRYB[4][16] ), .YS(\SUMB[4][16] ) );
  FAX1 S2_6_13 ( .A(n97), .B(\CARRYB[5][13] ), .C(\SUMB[5][14] ), .YC(
        \CARRYB[6][13] ), .YS(\SUMB[6][13] ) );
  FAX1 S2_5_14 ( .A(n98), .B(\CARRYB[4][14] ), .C(\SUMB[4][15] ), .YC(
        \CARRYB[5][14] ), .YS(\SUMB[5][14] ) );
  FAX1 S2_4_15 ( .A(n99), .B(\CARRYB[3][15] ), .C(\SUMB[3][16] ), .YC(
        \CARRYB[4][15] ), .YS(\SUMB[4][15] ) );
  FAX1 S2_3_16 ( .A(n102), .B(\CARRYB[2][16] ), .C(\SUMB[2][17] ), .YC(
        \CARRYB[3][16] ), .YS(\SUMB[3][16] ) );
  FAX1 S2_5_13 ( .A(n98), .B(\CARRYB[4][13] ), .C(\SUMB[4][14] ), .YC(
        \CARRYB[5][13] ), .YS(\SUMB[5][13] ) );
  FAX1 S2_4_14 ( .A(n99), .B(\CARRYB[3][14] ), .C(\SUMB[3][15] ), .YC(
        \CARRYB[4][14] ), .YS(\SUMB[4][14] ) );
  FAX1 S2_3_15 ( .A(n102), .B(\CARRYB[2][15] ), .C(\SUMB[2][16] ), .YC(
        \CARRYB[3][15] ), .YS(\SUMB[3][15] ) );
  FAX1 S2_2_16 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][16] ), .YS(
        \SUMB[2][16] ) );
  FAX1 S2_4_13 ( .A(n99), .B(\CARRYB[3][13] ), .C(\SUMB[3][14] ), .YC(
        \CARRYB[4][13] ), .YS(\SUMB[4][13] ) );
  FAX1 S2_3_14 ( .A(n102), .B(\CARRYB[2][14] ), .C(\SUMB[2][15] ), .YC(
        \CARRYB[3][14] ), .YS(\SUMB[3][14] ) );
  FAX1 S2_2_15 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][15] ), .YS(
        \SUMB[2][15] ) );
  FAX1 S2_3_13 ( .A(n102), .B(\CARRYB[2][13] ), .C(\SUMB[2][14] ), .YC(
        \CARRYB[3][13] ), .YS(\SUMB[3][13] ) );
  FAX1 S2_2_14 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][14] ), .YS(
        \SUMB[2][14] ) );
  FAX1 S2_2_13 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][13] ), .YS(
        \SUMB[2][13] ) );
  XOR2X1 U168 ( .A(\SUMB[7][18] ), .B(\CARRYB[7][17] ), .Y(\A1[23] ) );
  AND2X1 U52 ( .A(\CARRYB[7][17] ), .B(\SUMB[7][18] ), .Y(n31) );
  FAX1 S4_18 ( .A(n106), .B(\CARRYB[6][18] ), .C(\SUMB[6][19] ), .YC(
        \CARRYB[7][18] ), .YS(\SUMB[7][18] ) );
  FAX1 S2_6_19 ( .A(n97), .B(\CARRYB[5][19] ), .C(\SUMB[5][20] ), .YC(
        \CARRYB[6][19] ), .YS(\SUMB[6][19] ) );
  FAX1 S2_5_20 ( .A(n98), .B(\CARRYB[4][20] ), .C(\SUMB[4][21] ), .YC(
        \CARRYB[5][20] ), .YS(\SUMB[5][20] ) );
  FAX1 S4_17 ( .A(n106), .B(\CARRYB[6][17] ), .C(\SUMB[6][18] ), .YC(
        \CARRYB[7][17] ), .YS(\SUMB[7][17] ) );
  FAX1 S2_6_18 ( .A(n97), .B(\CARRYB[5][18] ), .C(\SUMB[5][19] ), .YC(
        \CARRYB[6][18] ), .YS(\SUMB[6][18] ) );
  FAX1 S2_5_19 ( .A(n98), .B(\CARRYB[4][19] ), .C(\SUMB[4][20] ), .YC(
        \CARRYB[5][19] ), .YS(\SUMB[5][19] ) );
  FAX1 S2_4_20 ( .A(n99), .B(\CARRYB[3][20] ), .C(\SUMB[3][21] ), .YC(
        \CARRYB[4][20] ), .YS(\SUMB[4][20] ) );
  FAX1 S2_6_17 ( .A(n97), .B(\CARRYB[5][17] ), .C(\SUMB[5][18] ), .YC(
        \CARRYB[6][17] ), .YS(\SUMB[6][17] ) );
  FAX1 S2_5_18 ( .A(n98), .B(\CARRYB[4][18] ), .C(\SUMB[4][19] ), .YC(
        \CARRYB[5][18] ), .YS(\SUMB[5][18] ) );
  FAX1 S2_4_19 ( .A(n99), .B(\CARRYB[3][19] ), .C(\SUMB[3][20] ), .YC(
        \CARRYB[4][19] ), .YS(\SUMB[4][19] ) );
  FAX1 S2_3_20 ( .A(n102), .B(\CARRYB[2][20] ), .C(\SUMB[2][21] ), .YC(
        \CARRYB[3][20] ), .YS(\SUMB[3][20] ) );
  FAX1 S2_5_17 ( .A(n98), .B(\CARRYB[4][17] ), .C(\SUMB[4][18] ), .YC(
        \CARRYB[5][17] ), .YS(\SUMB[5][17] ) );
  FAX1 S2_4_18 ( .A(n99), .B(\CARRYB[3][18] ), .C(\SUMB[3][19] ), .YC(
        \CARRYB[4][18] ), .YS(\SUMB[4][18] ) );
  FAX1 S2_3_19 ( .A(n102), .B(\CARRYB[2][19] ), .C(\SUMB[2][20] ), .YC(
        \CARRYB[3][19] ), .YS(\SUMB[3][19] ) );
  FAX1 S2_2_20 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][20] ), .YS(
        \SUMB[2][20] ) );
  FAX1 S2_4_17 ( .A(n99), .B(\CARRYB[3][17] ), .C(\SUMB[3][18] ), .YC(
        \CARRYB[4][17] ), .YS(\SUMB[4][17] ) );
  FAX1 S2_3_18 ( .A(n102), .B(\CARRYB[2][18] ), .C(\SUMB[2][19] ), .YC(
        \CARRYB[3][18] ), .YS(\SUMB[3][18] ) );
  FAX1 S2_2_19 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][19] ), .YS(
        \SUMB[2][19] ) );
  FAX1 S2_3_17 ( .A(n102), .B(\CARRYB[2][17] ), .C(\SUMB[2][18] ), .YC(
        \CARRYB[3][17] ), .YS(\SUMB[3][17] ) );
  FAX1 S2_2_18 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][18] ), .YS(
        \SUMB[2][18] ) );
  FAX1 S2_2_17 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][17] ), .YS(
        \SUMB[2][17] ) );
  XOR2X1 U164 ( .A(\SUMB[7][22] ), .B(\CARRYB[7][21] ), .Y(\A1[27] ) );
  AND2X1 U55 ( .A(\CARRYB[7][21] ), .B(\SUMB[7][22] ), .Y(n29) );
  FAX1 S4_22 ( .A(n106), .B(\CARRYB[6][22] ), .C(\SUMB[6][23] ), .YC(
        \CARRYB[7][22] ), .YS(\SUMB[7][22] ) );
  FAX1 S2_6_23 ( .A(n97), .B(\CARRYB[5][23] ), .C(\SUMB[5][24] ), .YC(
        \CARRYB[6][23] ), .YS(\SUMB[6][23] ) );
  FAX1 S2_5_24 ( .A(n98), .B(\CARRYB[4][24] ), .C(\SUMB[4][25] ), .YC(
        \CARRYB[5][24] ), .YS(\SUMB[5][24] ) );
  FAX1 S4_21 ( .A(n106), .B(\CARRYB[6][21] ), .C(\SUMB[6][22] ), .YC(
        \CARRYB[7][21] ), .YS(\SUMB[7][21] ) );
  FAX1 S2_6_22 ( .A(n97), .B(\CARRYB[5][22] ), .C(\SUMB[5][23] ), .YC(
        \CARRYB[6][22] ), .YS(\SUMB[6][22] ) );
  FAX1 S2_5_23 ( .A(n98), .B(\CARRYB[4][23] ), .C(\SUMB[4][24] ), .YC(
        \CARRYB[5][23] ), .YS(\SUMB[5][23] ) );
  FAX1 S2_4_24 ( .A(n99), .B(\CARRYB[3][24] ), .C(\SUMB[3][25] ), .YC(
        \CARRYB[4][24] ), .YS(\SUMB[4][24] ) );
  FAX1 S2_6_21 ( .A(n97), .B(\CARRYB[5][21] ), .C(\SUMB[5][22] ), .YC(
        \CARRYB[6][21] ), .YS(\SUMB[6][21] ) );
  FAX1 S2_5_22 ( .A(n98), .B(\CARRYB[4][22] ), .C(\SUMB[4][23] ), .YC(
        \CARRYB[5][22] ), .YS(\SUMB[5][22] ) );
  FAX1 S2_4_23 ( .A(n99), .B(\CARRYB[3][23] ), .C(\SUMB[3][24] ), .YC(
        \CARRYB[4][23] ), .YS(\SUMB[4][23] ) );
  FAX1 S2_3_24 ( .A(n102), .B(\CARRYB[2][24] ), .C(\SUMB[2][25] ), .YC(
        \CARRYB[3][24] ), .YS(\SUMB[3][24] ) );
  FAX1 S2_5_21 ( .A(n98), .B(\CARRYB[4][21] ), .C(\SUMB[4][22] ), .YC(
        \CARRYB[5][21] ), .YS(\SUMB[5][21] ) );
  FAX1 S2_4_22 ( .A(n99), .B(\CARRYB[3][22] ), .C(\SUMB[3][23] ), .YC(
        \CARRYB[4][22] ), .YS(\SUMB[4][22] ) );
  FAX1 S2_3_23 ( .A(n102), .B(\CARRYB[2][23] ), .C(\SUMB[2][24] ), .YC(
        \CARRYB[3][23] ), .YS(\SUMB[3][23] ) );
  FAX1 S2_2_24 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][24] ), .YS(
        \SUMB[2][24] ) );
  FAX1 S2_4_21 ( .A(n99), .B(\CARRYB[3][21] ), .C(\SUMB[3][22] ), .YC(
        \CARRYB[4][21] ), .YS(\SUMB[4][21] ) );
  FAX1 S2_3_22 ( .A(n102), .B(\CARRYB[2][22] ), .C(\SUMB[2][23] ), .YC(
        \CARRYB[3][22] ), .YS(\SUMB[3][22] ) );
  FAX1 S2_2_23 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][23] ), .YS(
        \SUMB[2][23] ) );
  FAX1 S2_3_21 ( .A(n102), .B(\CARRYB[2][21] ), .C(\SUMB[2][22] ), .YC(
        \CARRYB[3][21] ), .YS(\SUMB[3][21] ) );
  FAX1 S2_2_22 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][22] ), .YS(
        \SUMB[2][22] ) );
  FAX1 S2_2_21 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][21] ), .YS(
        \SUMB[2][21] ) );
  XOR2X1 U160 ( .A(\SUMB[7][26] ), .B(\CARRYB[7][25] ), .Y(\A1[31] ) );
  AND2X1 U36 ( .A(\CARRYB[7][25] ), .B(\SUMB[7][26] ), .Y(n8) );
  FAX1 S4_26 ( .A(n106), .B(\CARRYB[6][26] ), .C(\SUMB[6][27] ), .YC(
        \CARRYB[7][26] ), .YS(\SUMB[7][26] ) );
  FAX1 S2_6_27 ( .A(n97), .B(\CARRYB[5][27] ), .C(\SUMB[5][28] ), .YC(
        \CARRYB[6][27] ), .YS(\SUMB[6][27] ) );
  FAX1 S2_5_28 ( .A(n98), .B(\CARRYB[4][28] ), .C(\SUMB[4][29] ), .YC(
        \CARRYB[5][28] ), .YS(\SUMB[5][28] ) );
  FAX1 S4_25 ( .A(n106), .B(\CARRYB[6][25] ), .C(\SUMB[6][26] ), .YC(
        \CARRYB[7][25] ), .YS(\SUMB[7][25] ) );
  FAX1 S2_6_26 ( .A(n97), .B(\CARRYB[5][26] ), .C(\SUMB[5][27] ), .YC(
        \CARRYB[6][26] ), .YS(\SUMB[6][26] ) );
  FAX1 S2_5_27 ( .A(n98), .B(\CARRYB[4][27] ), .C(\SUMB[4][28] ), .YC(
        \CARRYB[5][27] ), .YS(\SUMB[5][27] ) );
  FAX1 S2_4_28 ( .A(n99), .B(\CARRYB[3][28] ), .C(\SUMB[3][29] ), .YC(
        \CARRYB[4][28] ), .YS(\SUMB[4][28] ) );
  FAX1 S2_6_25 ( .A(n97), .B(\CARRYB[5][25] ), .C(\SUMB[5][26] ), .YC(
        \CARRYB[6][25] ), .YS(\SUMB[6][25] ) );
  FAX1 S2_5_26 ( .A(n98), .B(\CARRYB[4][26] ), .C(\SUMB[4][27] ), .YC(
        \CARRYB[5][26] ), .YS(\SUMB[5][26] ) );
  FAX1 S2_4_27 ( .A(n99), .B(\CARRYB[3][27] ), .C(\SUMB[3][28] ), .YC(
        \CARRYB[4][27] ), .YS(\SUMB[4][27] ) );
  FAX1 S2_3_28 ( .A(n102), .B(\CARRYB[2][28] ), .C(\SUMB[2][29] ), .YC(
        \CARRYB[3][28] ), .YS(\SUMB[3][28] ) );
  FAX1 S2_5_25 ( .A(n98), .B(\CARRYB[4][25] ), .C(\SUMB[4][26] ), .YC(
        \CARRYB[5][25] ), .YS(\SUMB[5][25] ) );
  FAX1 S2_4_26 ( .A(n99), .B(\CARRYB[3][26] ), .C(\SUMB[3][27] ), .YC(
        \CARRYB[4][26] ), .YS(\SUMB[4][26] ) );
  FAX1 S2_3_27 ( .A(n102), .B(\CARRYB[2][27] ), .C(\SUMB[2][28] ), .YC(
        \CARRYB[3][27] ), .YS(\SUMB[3][27] ) );
  FAX1 S2_2_28 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][28] ), .YS(
        \SUMB[2][28] ) );
  FAX1 S2_4_25 ( .A(n99), .B(\CARRYB[3][25] ), .C(\SUMB[3][26] ), .YC(
        \CARRYB[4][25] ), .YS(\SUMB[4][25] ) );
  FAX1 S2_3_26 ( .A(n102), .B(\CARRYB[2][26] ), .C(\SUMB[2][27] ), .YC(
        \CARRYB[3][26] ), .YS(\SUMB[3][26] ) );
  FAX1 S2_2_27 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][27] ), .YS(
        \SUMB[2][27] ) );
  FAX1 S2_3_25 ( .A(n102), .B(\CARRYB[2][25] ), .C(\SUMB[2][26] ), .YC(
        \CARRYB[3][25] ), .YS(\SUMB[3][25] ) );
  FAX1 S2_2_26 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][26] ), .YS(
        \SUMB[2][26] ) );
  FAX1 S2_2_25 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][25] ), .YS(
        \SUMB[2][25] ) );
  XOR2X1 U156 ( .A(\SUMB[7][30] ), .B(\CARRYB[7][29] ), .Y(\A1[35] ) );
  AND2X1 U43 ( .A(\CARRYB[7][29] ), .B(\SUMB[7][30] ), .Y(n4) );
  FAX1 S5_30 ( .A(n106), .B(\CARRYB[6][30] ), .C(n97), .YC(\CARRYB[7][30] ), 
        .YS(\SUMB[7][30] ) );
  FAX1 S4_29 ( .A(n106), .B(\CARRYB[6][29] ), .C(\SUMB[6][30] ), .YC(
        \CARRYB[7][29] ), .YS(\SUMB[7][29] ) );
  FAX1 S3_6_30 ( .A(n97), .B(\CARRYB[5][30] ), .C(n98), .YC(\CARRYB[6][30] ), 
        .YS(\SUMB[6][30] ) );
  FAX1 S2_6_29 ( .A(n97), .B(\CARRYB[5][29] ), .C(\SUMB[5][30] ), .YC(
        \CARRYB[6][29] ), .YS(\SUMB[6][29] ) );
  FAX1 S3_5_30 ( .A(n98), .B(\CARRYB[4][30] ), .C(n99), .YC(\CARRYB[5][30] ), 
        .YS(\SUMB[5][30] ) );
  FAX1 S2_5_29 ( .A(n98), .B(\CARRYB[4][29] ), .C(\SUMB[4][30] ), .YC(
        \CARRYB[5][29] ), .YS(\SUMB[5][29] ) );
  FAX1 S3_4_30 ( .A(n99), .B(\CARRYB[3][30] ), .C(n102), .YC(\CARRYB[4][30] ), 
        .YS(\SUMB[4][30] ) );
  FAX1 S2_4_29 ( .A(n99), .B(\CARRYB[3][29] ), .C(\SUMB[3][30] ), .YC(
        \CARRYB[4][29] ), .YS(\SUMB[4][29] ) );
  FAX1 S3_3_30 ( .A(n102), .B(\CARRYB[2][30] ), .C(n103), .YC(\CARRYB[3][30] ), 
        .YS(\SUMB[3][30] ) );
  FAX1 S2_3_29 ( .A(n102), .B(\CARRYB[2][29] ), .C(\SUMB[2][30] ), .YC(
        \CARRYB[3][29] ), .YS(\SUMB[3][29] ) );
  FAX1 S3_2_30 ( .A(n103), .B(n105), .C(n145), .YC(\CARRYB[2][30] ), .YS(
        \SUMB[2][30] ) );
  FAX1 S2_2_29 ( .A(n103), .B(n105), .C(n101), .YC(\CARRYB[2][29] ), .YS(
        \SUMB[2][29] ) );
  NOR2X1 U145 ( .A(n109), .B(n107), .Y(n114) );
  AND2X1 U144 ( .A(A[1]), .B(B[9]), .Y(n145) );
  NOR2X1 U33 ( .A(n107), .B(n110), .Y(n143) );
  NOR2X1 U32 ( .A(n107), .B(n111), .Y(n142) );
  NOR2X1 U31 ( .A(n107), .B(n112), .Y(n141) );
  NOR2X1 U30 ( .A(n107), .B(n113), .Y(n140) );
  NOR2X1 U29 ( .A(n107), .B(n144), .Y(n139) );
  NOR2X1 U155 ( .A(n107), .B(n146), .Y(n138) );
  BUFX4 U12 ( .A(n139), .Y(n97) );
  BUFX4 U13 ( .A(n140), .Y(n98) );
  BUFX4 U14 ( .A(n141), .Y(n99) );
  XOR2X1 U15 ( .A(n108), .B(n145), .Y(n100) );
  INVX2 U16 ( .A(n100), .Y(n101) );
  BUFX4 U17 ( .A(n142), .Y(n102) );
  BUFX4 U18 ( .A(n143), .Y(n103) );
  NAND2X1 U19 ( .A(n145), .B(n114), .Y(n104) );
  INVX4 U20 ( .A(n104), .Y(n105) );
  BUFX4 U21 ( .A(n138), .Y(n106) );
  INVX2 U22 ( .A(B[9]), .Y(n107) );
  INVX2 U23 ( .A(n114), .Y(n108) );
  INVX2 U24 ( .A(A[0]), .Y(n109) );
  INVX2 U25 ( .A(A[2]), .Y(n110) );
  INVX2 U26 ( .A(A[3]), .Y(n111) );
  INVX2 U27 ( .A(A[4]), .Y(n112) );
  INVX2 U28 ( .A(A[5]), .Y(n113) );
  INVX2 U34 ( .A(A[6]), .Y(n144) );
  INVX2 U143 ( .A(A[7]), .Y(n146) );
  INVX2 U182 ( .A(B[0]), .Y(n147) );
  INVX2 U183 ( .A(B[1]), .Y(n148) );
  INVX2 U184 ( .A(B[2]), .Y(n149) );
  INVX2 U185 ( .A(B[3]), .Y(n150) );
  INVX2 U186 ( .A(B[4]), .Y(n151) );
  INVX2 U187 ( .A(B[5]), .Y(n152) );
  INVX2 U188 ( .A(B[6]), .Y(n153) );
  INVX2 U189 ( .A(B[7]), .Y(n154) );
endmodule


module CannyEdge ( dAddrRegRow, dAddrRegCol, bWE, bCE, InData, OutData, OPMode, 
        bOPEnable, dReadReg, dWriteReg, clk, rst_b );
  input [2:0] dAddrRegRow;
  input [2:0] dAddrRegCol;
  input [7:0] InData;
  output [7:0] OutData;
  input [2:0] OPMode;
  input [3:0] dReadReg;
  input [3:0] dWriteReg;
  input bWE, bCE, bOPEnable, clk, rst_b;
  wire   \regX[0][7] , \regX[0][6] , \regX[0][5] , \regX[0][4] , \regX[0][3] ,
         \regX[0][2] , \regX[0][1] , \regX[0][0] , \regX[1][7] , \regX[1][6] ,
         \regX[1][5] , \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] ,
         \regX[1][0] , \regX[3][7] , \regX[3][6] , \regX[3][5] , \regX[3][4] ,
         \regX[3][3] , \regX[3][2] , \regX[3][1] , \regX[3][0] , \regX[5][7] ,
         \regX[5][6] , \regX[5][5] , \regX[5][4] , \regX[5][3] , \regX[5][2] ,
         \regX[5][1] , \regX[5][0] , \regX[6][7] , \regX[6][6] , \regX[6][5] ,
         \regX[6][4] , \regX[6][3] , \regX[6][2] , \regX[6][1] , \regX[6][0] ,
         \regX[7][7] , \regX[7][6] , \regX[7][5] , \regX[7][4] , \regX[7][3] ,
         \regX[7][2] , \regX[7][1] , \regX[7][0] , \regX[8][7] , \regX[8][6] ,
         \regX[8][5] , \regX[8][4] , \regX[8][3] , \regX[8][2] , \regX[8][1] ,
         \regX[8][0] , \regX[9][7] , \regX[9][6] , \regX[9][5] , \regX[9][4] ,
         \regX[9][3] , \regX[9][2] , \regX[9][1] , \regX[9][0] , \regX[11][7] ,
         \regX[11][6] , \regX[11][5] , \regX[11][4] , \regX[11][3] ,
         \regX[11][2] , \regX[11][1] , \regX[11][0] , \regX[13][7] ,
         \regX[13][6] , \regX[13][5] , \regX[13][4] , \regX[13][3] ,
         \regX[13][2] , \regX[13][1] , \regX[13][0] , \regX[15][7] ,
         \regX[15][6] , \regX[15][5] , \regX[15][4] , \regX[15][3] ,
         \regX[15][2] , \regX[15][1] , \regX[15][0] , \regX[16][7] ,
         \regX[16][6] , \regX[16][5] , \regX[16][4] , \regX[16][3] ,
         \regX[16][2] , \regX[16][1] , \regX[16][0] , \regX[17][7] ,
         \regX[17][6] , \regX[17][5] , \regX[17][4] , \regX[17][3] ,
         \regX[17][2] , \regX[17][1] , \regX[17][0] , \regX[18][7] ,
         \regX[18][6] , \regX[18][5] , \regX[18][4] , \regX[18][3] ,
         \regX[18][2] , \regX[18][1] , \regX[18][0] , \regX[19][7] ,
         \regX[19][6] , \regX[19][5] , \regX[19][4] , \regX[19][3] ,
         \regX[19][2] , \regX[19][1] , \regX[19][0] , \regX[20][7] ,
         \regX[20][6] , \regX[20][5] , \regX[20][4] , \regX[20][3] ,
         \regX[20][2] , \regX[20][1] , \regX[20][0] , \regX[21][7] ,
         \regX[21][6] , \regX[21][5] , \regX[21][4] , \regX[21][3] ,
         \regX[21][2] , \regX[21][1] , \regX[21][0] , \regX[22][7] ,
         \regX[22][6] , \regX[22][5] , \regX[22][4] , \regX[22][3] ,
         \regX[22][2] , \regX[22][1] , \regX[22][0] , \regX[23][7] ,
         \regX[23][6] , \regX[23][5] , \regX[23][4] , \regX[23][3] ,
         \regX[23][2] , \regX[23][1] , \regX[23][0] , \regX[24][7] ,
         \regX[24][6] , \regX[24][5] , \regX[24][4] , \regX[24][3] ,
         \regX[24][2] , \regX[24][1] , \regX[24][0] , \regY[6][7] ,
         \regY[6][6] , \regY[6][5] , \regY[6][4] , \regY[6][3] , \regY[6][2] ,
         \regY[6][1] , \regY[6][0] , N971, N972, N973, N974, N975, N976, N977,
         N978, N979, N980, N981, N982, N983, \Out_bThres[0] , N1343, N1344,
         N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354,
         N1355, N1356, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382,
         N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397,
         N1398, N1399, N1400, N1401, N1402, N1408, N1409, N1410, N1411, N1412,
         N1413, N1414, N1415, N1416, N1417, N1433, N1434, N1435, N1436, N1437,
         N1438, N1439, N1440, N1510, N1511, N1512, N1513, N1514, N1515, N1516,
         N1517, N1518, N1519, N1520, N1521, N1522, N1542, N1543, N1544, N1545,
         N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1570, N1571, N1572,
         N1573, N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582,
         N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1645, N1646,
         N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656,
         N1677, N1678, N1679, N1680, N1681, N1682, N1683, N1684, N1707, N1708,
         N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1735, N1736,
         N1737, N1738, N1739, N1740, N1741, N1742, N1765, N1766, N1767, N1768,
         N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N2048, N2049,
         N2050, N2051, N2052, N2053, N2054, N2055, N2091, N2092, N2093, N2094,
         N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104,
         N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114,
         N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2155, N2156,
         N2157, N2158, N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166,
         N2167, N2168, N2169, N2170, N2171, N2236, N2237, N2238, N2239, N2240,
         N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250,
         N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260,
         N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270,
         N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280,
         N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290,
         N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300,
         N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310,
         N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320,
         N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330,
         N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340,
         N2341, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393,
         N2394, N2395, N2396, N2397, N2398, N2399, N2513, N2514, N2515, N2516,
         N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526,
         N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536,
         N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2549, N2558,
         N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568,
         N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2648, N2746,
         N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756,
         N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766,
         N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776,
         N2777, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832,
         N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2874,
         N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889,
         N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899,
         N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909,
         N2910, N2911, N2945, N3089, N3090, N3091, N3092, N3093, N3189, N3190,
         N3191, N3192, N3193, N3194, N3336, N3340, N3341, N3342, N3343, N3359,
         N3441, N3442, N3443, N3772, N3773, N3775, N3776, N3778, N3779, N3781,
         N3782, N3784, N3785, N3787, N3788, N3790, N3791, N3793, N3794, N3796,
         N3797, N3799, N3800, N3802, N3803, N3805, N3806, N3808, N3809, N3811,
         N3812, N3814, N3815, N3817, N3818, N3820, N3821, N3823, N3824, N3826,
         N3827, N3829, N3830, N3832, N3833, N3835, N3836, N3838, N3839, N3841,
         N3842, N3844, N3845, N3847, N3848, N3850, N3851, N3853, N3854, N3856,
         N3857, N3859, N3860, N3862, N3863, N3865, N3866, N3868, N3869, N3871,
         N3872, N3874, N3875, N3877, N3878, N3880, N3881, N3883, N3884, N3886,
         N3887, N3889, N3890, N3892, N3893, N3895, N3896, N3898, N3899, N3901,
         N3902, N3904, N3905, N3907, N3908, N3910, N3911, N3913, N3914, N3916,
         N3917, N3919, N3920, N3922, N3923, N3925, N3926, N3928, N3929, N3931,
         N3932, N3934, N3935, N3937, N3938, N3940, N3941, N3943, N3944, N3946,
         N3947, N3949, N3950, N3952, N3953, N3955, N3956, N3958, N3959, N3961,
         N3962, N3964, N3965, N3967, N3968, N3970, N3971, N3973, N3974, N3976,
         N3977, N3979, N3980, N3982, N3983, N3985, N3986, N3988, N3989, N3991,
         N3992, N3994, N3995, N3997, N3998, N4000, N4001, N4003, N4004, N4006,
         N4007, N4009, N4010, N4012, N4013, N4015, N4016, N4018, N4019, N4021,
         N4022, N4024, N4025, N4027, N4028, N4030, N4031, N4033, N4034, N4036,
         N4037, N4039, N4040, N4042, N4043, N4045, N4046, N4048, N4049, N4051,
         N4052, N4054, N4055, N4057, N4058, N4060, N4061, N4063, N4064, N4066,
         N4067, N4069, N4070, N4072, N4073, N4075, N4076, N4078, N4079, N4081,
         N4082, N4084, N4085, N4087, N4088, N4090, N4091, N4093, N4094, N4096,
         N4097, N4099, N4100, N4102, N4103, N4105, N4106, N4108, N4109, N4111,
         N4112, N4114, N4115, N4117, N4118, N4120, N4121, N4123, N4124, N4126,
         N4127, N4129, N4130, N4132, N4133, N4135, N4136, N4138, N4139, N4141,
         N4142, N4144, N4145, N4147, N4148, N4150, N4151, N4153, N4154, N4156,
         N4157, N4159, N4160, N4162, N4163, N4165, N4166, N4168, N4169, N4171,
         N4172, N4174, N4175, N4177, N4178, N4180, N4181, N4183, N4184, N4186,
         N4187, N4189, N4190, N4192, N4193, N4195, N4196, N4198, N4199, N4201,
         N4202, N4204, N4205, N4207, N4208, N4210, N4211, N4213, N4214, N4216,
         N4217, N4219, N4220, N4222, N4223, N4225, N4226, N4228, N4229, N4231,
         N4232, N4234, N4235, N4237, N4238, N4240, N4241, N4243, N4244, N4246,
         N4247, N4249, N4250, N4252, N4253, N4255, N4256, N4258, N4259, N4261,
         N4262, N4264, N4265, N4267, N4268, N4270, N4271, N4273, N4274, N4276,
         N4277, N4279, N4280, N4282, N4283, N4285, N4286, N4288, N4289, N4291,
         N4292, N4294, N4295, N4297, N4298, N4300, N4301, N4303, N4304, N4306,
         N4307, N4309, N4310, N4312, N4313, N4315, N4316, N4318, N4319, N4321,
         N4322, N4324, N4325, N4327, N4328, N4330, N4331, N4333, N4334, N4336,
         N4337, N4339, N4340, N4342, N4343, N4345, N4346, N4348, N4349, N4351,
         N4352, N4354, N4355, N4357, N4358, N4360, N4361, N4363, N4364, N4366,
         N4367, N4369, N4370, N4372, N4373, N4375, N4376, N4378, N4379, N4381,
         N4382, N4384, N4385, N4387, N4388, N4390, N4391, N4393, N4394, N4396,
         N4397, N4399, N4400, N4402, N4403, N4405, N4406, N4408, N4409, N4411,
         N4412, N4414, N4415, N4417, N4418, N4420, N4421, N4423, N4424, N4426,
         N4427, N4429, N4430, N4432, N4433, N4435, N4436, N4438, N4439, N4441,
         N4442, N4444, N4445, N4447, N4448, N4450, N4451, N4453, N4454, N4456,
         N4457, N4459, N4460, N4462, N4463, N4465, N4466, N4468, N4469, N4471,
         N4472, N4474, N4475, N4477, N4478, N4480, N4481, N4483, N4484, N4486,
         N4487, N4489, N4490, N4495, N4496, N4501, N4502, \U3/U63/Z_0 ,
         \U3/U63/Z_1 , \U3/U63/Z_2 , \U3/U63/Z_3 , \U3/U63/Z_4 , \U3/U63/Z_5 ,
         \U3/U63/Z_6 , \U3/U63/Z_7 , \U3/U64/Z_0 , \U3/U64/Z_1 , \U3/U64/Z_2 ,
         \U3/U64/Z_3 , \U3/U64/Z_4 , \U3/U64/Z_5 , \U3/U64/Z_6 , \U3/U64/Z_7 ,
         \U3/U65/Z_0 , \U3/U65/Z_1 , \U3/U65/Z_2 , \U3/U65/Z_3 , \U3/U65/Z_4 ,
         \U3/U65/Z_5 , \U3/U65/Z_6 , \U3/U65/Z_7 , \U3/U68/Z_15 ,
         \U3/U68/Z_16 , \U3/U68/Z_17 , \U3/U68/Z_18 , \U3/U68/Z_19 ,
         \U3/U68/Z_20 , \U3/U68/Z_21 , \U3/U68/Z_22 , \U3/U68/Z_23 ,
         \U3/U68/Z_24 , \U3/U68/Z_25 , \U3/U68/Z_26 , \U3/U68/Z_27 ,
         \U3/U68/Z_28 , \U3/U68/Z_29 , \U3/U68/Z_30 , \U3/U68/Z_31 ,
         \U3/U69/Z_0 , \U3/U69/Z_1 , \U3/U69/Z_2 , \U3/U69/Z_3 , \U3/U69/Z_4 ,
         \U3/U69/Z_5 , \U3/U69/Z_6 , \U3/U69/Z_7 , \U3/U69/Z_8 , \U3/U69/Z_9 ,
         \U3/U69/Z_10 , \U3/U69/Z_11 , \U3/U69/Z_12 , \U3/U69/Z_13 ,
         \U3/U70/Z_0 , \U3/U70/Z_1 , \U3/U70/Z_2 , \U3/U70/Z_3 , \U3/U70/Z_4 ,
         \U3/U70/Z_5 , \U3/U70/Z_6 , \U3/U70/Z_7 , \U3/U70/Z_8 , \U3/U71/Z_15 ,
         \U3/U71/Z_16 , \U3/U71/Z_17 , \U3/U71/Z_18 , \U3/U71/Z_19 ,
         \U3/U71/Z_20 , \U3/U71/Z_21 , \U3/U71/Z_22 , \U3/U71/Z_23 ,
         \U3/U71/Z_24 , \U3/U71/Z_25 , \U3/U71/Z_26 , \U3/U71/Z_27 ,
         \U3/U71/Z_28 , \U3/U71/Z_29 , \U3/U71/Z_30 , \U3/U71/Z_31 ,
         \U3/U72/Z_15 , \U3/U72/Z_16 , \U3/U72/Z_17 , \U3/U72/Z_18 ,
         \U3/U72/Z_19 , \U3/U72/Z_20 , \U3/U72/Z_21 , \U3/U72/Z_22 ,
         \U3/U72/Z_23 , \U3/U72/Z_24 , \U3/U72/Z_25 , \U3/U72/Z_26 ,
         \U3/U72/Z_27 , \U3/U72/Z_28 , \U3/U72/Z_29 , \U3/U72/Z_30 ,
         \U3/U72/Z_31 , \U3/U73/Z_15 , \U3/U73/Z_16 , \U3/U73/Z_17 ,
         \U3/U73/Z_18 , \U3/U73/Z_19 , \U3/U73/Z_20 , \U3/U73/Z_21 ,
         \U3/U73/Z_22 , \U3/U73/Z_23 , \U3/U73/Z_24 , \U3/U73/Z_25 ,
         \U3/U73/Z_26 , \U3/U73/Z_27 , \U3/U73/Z_28 , \U3/U73/Z_29 ,
         \U3/U73/Z_30 , \U3/U73/Z_31 , \U3/U74/Z_15 , \U3/U74/Z_16 ,
         \U3/U74/Z_17 , \U3/U74/Z_18 , \U3/U74/Z_19 , \U3/U74/Z_20 ,
         \U3/U74/Z_21 , \U3/U74/Z_22 , \U3/U74/Z_23 , \U3/U74/Z_24 ,
         \U3/U74/Z_25 , \U3/U74/Z_26 , \U3/U74/Z_27 , \U3/U74/Z_28 ,
         \U3/U74/Z_29 , \U3/U74/Z_30 , \U3/U74/Z_31 , \U3/U75/Z_0 ,
         \U3/U75/Z_1 , \U3/U75/Z_2 , \U3/U75/Z_3 , \U3/U75/Z_4 , \U3/U75/Z_5 ,
         \U3/U75/Z_6 , \U3/U75/Z_7 , \U3/U75/Z_8 , \U3/U75/Z_9 , \U3/U75/Z_10 ,
         \U3/U75/Z_11 , \U3/U75/Z_12 , \U3/U75/Z_13 , \U3/U75/Z_14 ,
         \U3/U76/Z_10 , \U3/U76/Z_11 , \U3/U76/Z_12 , \U3/U76/Z_13 ,
         \U3/U76/Z_14 , \U3/U77/Z_15 , \U3/U77/Z_16 , \U3/U77/Z_17 ,
         \U3/U77/Z_18 , \U3/U77/Z_19 , \U3/U77/Z_20 , \U3/U77/Z_21 ,
         \U3/U77/Z_22 , \U3/U77/Z_23 , \U3/U77/Z_24 , \U3/U77/Z_25 ,
         \U3/U77/Z_26 , \U3/U77/Z_27 , \U3/U77/Z_28 , \U3/U77/Z_29 ,
         \U3/U77/Z_30 , \U3/U77/Z_31 , \U3/U77/DATA2_15 , \U3/U77/DATA2_16 ,
         \U3/U77/DATA2_17 , \U3/U77/DATA2_18 , \U3/U77/DATA2_19 ,
         \U3/U77/DATA2_20 , \U3/U77/DATA2_21 , \U3/U77/DATA2_22 ,
         \U3/U77/DATA2_23 , \U3/U77/DATA2_24 , \U3/U77/DATA2_25 ,
         \U3/U77/DATA2_26 , \U3/U77/DATA2_27 , \U3/U77/DATA2_28 ,
         \U3/U77/DATA2_29 , \U3/U77/DATA2_30 , \U3/U77/DATA2_31 , \U3/U78/Z_0 ,
         \U3/U78/Z_1 , \U3/U78/Z_2 , \U3/U78/Z_3 , \U3/U78/Z_4 , \U3/U78/Z_5 ,
         \U3/U78/Z_6 , \U3/U78/Z_7 , \U3/U78/Z_8 , \U3/U78/Z_9 , \U3/U78/Z_10 ,
         \U3/U78/Z_11 , \U3/U78/Z_12 , \U3/U78/Z_13 , \U3/U78/Z_14 ,
         \U3/U78/Z_15 , \U3/U78/Z_16 , \U3/U78/Z_17 , \U3/U78/Z_18 ,
         \U3/U78/Z_19 , \U3/U78/Z_20 , \U3/U78/Z_21 , \U3/U78/Z_22 ,
         \U3/U78/Z_23 , \U3/U78/Z_24 , \U3/U78/Z_25 , \U3/U78/Z_26 ,
         \U3/U78/Z_27 , \U3/U78/Z_28 , \U3/U78/Z_29 , \U3/U78/Z_30 ,
         \U3/U78/Z_31 , \U3/U79/Z_0 , \U3/U79/Z_1 , \U3/U79/Z_2 , \U3/U79/Z_3 ,
         \U3/U79/Z_4 , \U3/U79/Z_5 , \U3/U79/Z_6 , \U3/U79/Z_7 , \U3/U79/Z_8 ,
         \U3/U79/Z_9 , \U3/U79/Z_10 , \U3/U79/Z_11 , \U3/U79/Z_12 ,
         \U3/U79/Z_13 , \U3/U79/Z_14 , \U3/U79/Z_15 , \U3/U79/Z_16 ,
         \U3/U79/Z_17 , \U3/U79/Z_18 , \U3/U79/Z_19 , \U3/U79/Z_20 ,
         \U3/U79/Z_21 , \U3/U79/Z_22 , \U3/U79/Z_23 , \U3/U79/Z_24 ,
         \U3/U79/Z_25 , \U3/U79/Z_26 , \U3/U79/Z_27 , \U3/U79/Z_28 ,
         \U3/U79/Z_29 , \U3/U79/Z_30 , \U3/U79/Z_31 , \U3/U81/Z_0 ,
         \U3/U81/Z_1 , \U3/U81/Z_2 , \U3/U81/Z_3 , \U3/U81/Z_4 , \U3/U81/Z_5 ,
         \U3/U81/Z_6 , \U3/U81/Z_7 , \U3/U82/Z_0 , \U3/U82/Z_1 , \U3/U82/Z_2 ,
         \U3/U82/Z_3 , \U3/U82/Z_4 , \U3/U82/Z_5 , \U3/U82/Z_6 , \U3/U82/Z_7 ,
         \U3/U82/Z_8 , \U3/U82/Z_9 , \U3/U82/Z_10 , \U3/U82/Z_11 ,
         \U3/U82/Z_12 , \U3/U82/Z_13 , \U3/U82/Z_14 , \U3/U82/Z_15 ,
         \U3/U82/Z_16 , \U3/U82/Z_17 , \U3/U82/Z_18 , \U3/U82/Z_19 ,
         \U3/U82/Z_20 , \U3/U82/Z_21 , \U3/U82/Z_22 , \U3/U82/Z_23 ,
         \U3/U82/Z_24 , \U3/U82/Z_25 , \U3/U82/Z_26 , \U3/U82/Z_27 ,
         \U3/U82/Z_28 , \U3/U82/Z_29 , \U3/U82/Z_30 , \U3/U82/Z_31 ,
         \U3/U84/Z_0 , \U3/U84/Z_1 , \U3/U84/Z_2 , \U3/U84/Z_3 , \U3/U84/Z_4 ,
         \U3/U84/Z_5 , \U3/U84/Z_6 , \U3/U84/Z_7 , \U3/U85/Z_0 , \U3/U85/Z_1 ,
         \U3/U85/Z_2 , \U3/U85/Z_3 , \U3/U85/Z_4 , \U3/U85/Z_5 , \U3/U85/Z_6 ,
         \U3/U85/Z_7 , \U3/U85/Z_8 , \U3/U85/Z_9 , \U3/U85/Z_10 ,
         \U3/U85/Z_11 , \U3/U85/Z_12 , \U3/U85/Z_13 , \U3/U85/Z_14 ,
         \U3/U85/Z_15 , \U3/U85/Z_16 , \U3/U85/Z_17 , \U3/U85/Z_18 ,
         \U3/U85/Z_19 , \U3/U85/Z_20 , \U3/U85/Z_21 , \U3/U85/Z_22 ,
         \U3/U85/Z_23 , \U3/U85/Z_24 , \U3/U85/Z_25 , \U3/U85/Z_26 ,
         \U3/U85/Z_27 , \U3/U85/Z_28 , \U3/U85/Z_29 , \U3/U85/Z_30 ,
         \U3/U85/Z_31 , \U3/U87/Z_0 , \U3/U87/Z_1 , \U3/U87/Z_2 , \U3/U87/Z_3 ,
         \U3/U87/Z_4 , \U3/U87/Z_5 , \U3/U87/Z_6 , \U3/U87/Z_7 , \U3/U88/Z_0 ,
         \U3/U88/Z_1 , \U3/U88/Z_2 , \U3/U88/Z_3 , \U3/U88/Z_4 , \U3/U88/Z_5 ,
         \U3/U88/Z_6 , \U3/U88/Z_7 , \U3/U88/Z_8 , \U3/U88/Z_9 , \U3/U88/Z_10 ,
         \U3/U88/Z_11 , \U3/U88/Z_12 , \U3/U88/Z_13 , \U3/U88/Z_14 ,
         \U3/U88/Z_15 , \U3/U88/Z_16 , \U3/U88/Z_17 , \U3/U88/Z_18 ,
         \U3/U88/Z_19 , \U3/U88/Z_20 , \U3/U88/Z_21 , \U3/U88/Z_22 ,
         \U3/U88/Z_23 , \U3/U88/Z_24 , \U3/U88/Z_25 , \U3/U88/Z_26 ,
         \U3/U88/Z_27 , \U3/U88/Z_28 , \U3/U88/Z_29 , \U3/U88/Z_30 ,
         \U3/U90/Z_0 , \U3/U91/Z_0 , \U3/U91/Z_1 , \U3/U91/Z_2 , \U3/U91/Z_3 ,
         \U3/U91/Z_4 , \U3/U91/Z_5 , \U3/U91/Z_6 , \U3/U91/Z_7 , \U3/U93/Z_0 ,
         \U3/U93/Z_1 , \U3/U93/Z_2 , \U3/U93/Z_3 , \U3/U93/Z_4 , \U3/U93/Z_5 ,
         \U3/U93/Z_6 , \U3/U93/Z_7 , \U3/U93/Z_8 , \U3/U93/Z_9 , \U3/U93/Z_10 ,
         \U3/U93/Z_11 , \U3/U93/Z_12 , \U3/U93/Z_13 , \U3/U93/Z_14 ,
         \U3/U93/Z_15 , \U3/U93/Z_16 , \U3/U93/Z_17 , \U3/U93/Z_18 ,
         \U3/U93/Z_19 , \U3/U93/Z_20 , \U3/U93/Z_21 , \U3/U93/Z_22 ,
         \U3/U93/Z_23 , \U3/U93/Z_24 , \U3/U93/Z_25 , \U3/U93/Z_26 ,
         \U3/U93/Z_27 , \U3/U93/Z_28 , \U3/U93/Z_29 , \U3/U93/Z_30 ,
         \U3/U93/Z_31 , \U3/U94/Z_0 , \U3/U94/Z_1 , \U3/U94/Z_2 , \U3/U94/Z_3 ,
         \U3/U94/Z_4 , \U3/U94/Z_5 , \U3/U94/Z_6 , \U3/U94/Z_7 , \U3/U94/Z_8 ,
         \U3/U94/Z_9 , \U3/U94/Z_10 , \U3/U94/Z_11 , \U3/U94/Z_12 ,
         \U3/U94/Z_13 , \U3/U94/Z_14 , \U3/U94/Z_15 , \U3/U94/Z_16 ,
         \U3/U94/Z_17 , \U3/U94/Z_18 , \U3/U94/Z_19 , \U3/U94/Z_20 ,
         \U3/U94/Z_21 , \U3/U94/Z_22 , \U3/U94/Z_23 , \U3/U94/Z_24 ,
         \U3/U94/Z_25 , \U3/U94/Z_26 , \U3/U94/Z_27 , \U3/U94/Z_28 ,
         \U3/U94/Z_29 , \U3/U94/Z_31 , \U3/U95/Z_0 , \U3/U96/Z_0 ,
         \U3/U97/Z_0 , \U3/U98/Z_0 , \U3/U98/Z_1 , \U3/U98/Z_2 , \U3/U98/Z_3 ,
         \U3/U98/Z_4 , \U3/U98/Z_5 , \U3/U98/Z_6 , \U3/U98/Z_7 , \U3/U100/Z_6 ,
         \U3/U101/Z_0 , \U3/U101/Z_3 , \U3/U101/Z_6 , \U3/U105/Z_0 ,
         \U3/U105/Z_1 , \U3/U105/Z_2 , \U3/U105/Z_3 , \U3/U106/Z_1 ,
         \U3/U106/Z_3 , \U3/U109/Z_2 , \U3/U110/Z_0 , \U3/U110/Z_1 ,
         \U3/U110/Z_2 , \U3/U110/Z_3 , \U3/U110/Z_4 , \U3/U110/Z_5 ,
         \U3/U110/Z_6 , \U3/U110/Z_7 , \U3/U118/Z_0 , \U3/U118/Z_1 ,
         \U3/U118/Z_2 , \U3/U118/Z_3 , \U3/U118/Z_4 , \U3/U118/Z_5 ,
         \U3/U118/Z_6 , \U3/U118/Z_7 , \U3/U118/Z_8 , \U3/U118/Z_9 ,
         \U3/U118/Z_10 , \U3/U118/Z_11 , \U3/U118/Z_12 , \U3/U118/Z_13 ,
         \U3/U118/Z_14 , \U3/U118/Z_15 , \U3/U118/Z_16 , \U3/U118/Z_17 ,
         \U3/U118/Z_18 , \U3/U118/Z_19 , \U3/U118/Z_20 , \U3/U118/Z_21 ,
         \U3/U118/Z_22 , \U3/U118/Z_23 , \U3/U118/Z_24 , \U3/U118/Z_25 ,
         \U3/U118/Z_26 , \U3/U118/Z_27 , \U3/U118/Z_28 , \U3/U118/Z_29 ,
         \U3/U118/Z_30 , \U3/U118/Z_31 , \U3/U119/Z_0 , \U3/U119/Z_1 ,
         \U3/U119/Z_2 , \U3/U119/Z_3 , \U3/U119/Z_4 , \U3/U119/Z_5 ,
         \U3/U119/Z_6 , \U3/U119/Z_7 , \U3/U119/Z_8 , \U3/U119/Z_9 ,
         \U3/U119/Z_10 , \U3/U119/Z_11 , \U3/U119/Z_12 , \U3/U119/Z_13 ,
         \U3/U119/Z_14 , \U3/U119/Z_15 , \U3/U119/Z_16 , \U3/U119/Z_17 ,
         \U3/U119/Z_18 , \U3/U119/Z_19 , \U3/U119/Z_20 , \U3/U119/Z_21 ,
         \U3/U119/Z_22 , \U3/U119/Z_23 , \U3/U119/Z_24 , \U3/U119/Z_25 ,
         \U3/U119/Z_26 , \U3/U119/Z_27 , \U3/U119/Z_28 , \U3/U119/Z_29 ,
         \U3/U119/Z_31 , \U3/U121/Z_0 , \U3/U121/Z_1 , \U3/U121/Z_2 ,
         \U3/U121/Z_3 , \U3/U121/Z_4 , \U3/U121/Z_5 , \U3/U121/Z_6 ,
         \U3/U121/Z_7 , \U3/U122/Z_0 , \U3/U122/Z_1 , \U3/U122/Z_2 ,
         \U3/U122/Z_3 , \U3/U122/Z_4 , \U3/U122/Z_5 , \U3/U122/Z_6 ,
         \U3/U122/Z_7 , \U3/U122/Z_8 , \U3/U122/Z_9 , \U3/U122/Z_10 ,
         \U3/U122/Z_11 , \U3/U122/Z_12 , \U3/U122/Z_13 , \U3/U122/Z_14 ,
         \U3/U122/Z_15 , \U3/U122/Z_16 , \U3/U122/Z_17 , \U3/U122/Z_18 ,
         \U3/U122/Z_19 , \U3/U122/Z_20 , \U3/U122/Z_21 , \U3/U122/Z_22 ,
         \U3/U122/Z_23 , \U3/U122/Z_24 , \U3/U122/Z_25 , \U3/U122/Z_26 ,
         \U3/U122/Z_27 , \U3/U122/Z_28 , \U3/U122/Z_29 , \U3/U124/Z_0 ,
         \U3/U125/Z_0 , \U3/U125/Z_1 , \U3/U125/Z_2 , \U3/U125/Z_3 ,
         \U3/U125/Z_4 , \U3/U125/Z_5 , \U3/U125/Z_6 , \U3/U125/Z_7 ,
         \U3/U134/Z_0 , \U3/U134/Z_1 , \U3/U134/Z_2 , \U3/U134/Z_3 ,
         \U3/U134/Z_4 , \U3/U134/Z_5 , \U3/U134/Z_6 , \U3/U134/Z_7 ,
         \U3/U134/Z_8 , \U3/U134/Z_9 , \U3/U134/Z_10 , \U3/U136/Z_0 , n4572,
         n4573, n4574, n4612, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n2980,
         N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814,
         N2813, N2812, N2811, N2810, N2481, N2480, N2479, N2478, N2477, N2476,
         N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466,
         N2465, N2464, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410,
         N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400,
         N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194,
         N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184,
         N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174,
         N2173, N2172, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147,
         N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137,
         N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127,
         N2126, N2125, N2124, N2123, N2090, N2089, N2088, N2087, N2086, N2085,
         N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2032,
         N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022,
         N2021, N2020, N2019, N2018, N2002, N2001, N2000, N1999, N1998, N1997,
         N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1972,
         N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962,
         N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952,
         N1951, N1950, N1949, N1942, N1941, N1940, N1939, N1938, N1937, N1936,
         N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926,
         N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1912, N1911,
         N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901,
         N1900, N1899, N1898, N1896, N1895, N1894, N1893, N1892, N1891, N1890,
         N1889, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874,
         N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864,
         N1863, N1862, N1861, N1860, N1859, N1858, N1852, N1851, N1850, N1849,
         N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839,
         N1838, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828,
         N1827, N1826, N1825, N1824, N1822, N1821, N1820, N1819, N1818, N1817,
         N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1806, N1805,
         N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795,
         N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785,
         N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1762, N1761, N1760,
         N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750,
         N1749, N1748, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725,
         N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1672, N1671, N1670,
         N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660,
         N1659, N1658, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635,
         N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1612, N1611, N1610,
         N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600,
         N1599, N1598, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589,
         N1588, N1587, N1586, N1585, N1584, N1583, N1569, N1568, N1566, N1565,
         N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555,
         N1554, N1553, N1541, N1540, N1539, N1536, N1535, N1534, N1533, N1532,
         N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1509, N1506,
         N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496,
         N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486,
         N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1462, N1461,
         N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451,
         N1450, N1449, N1448, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3740, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n5089, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737;
  wire   [7:0] Out_gf;
  wire   [1:0] IntSignal;
  wire   [14:7] tpSum;
  wire   [31:0] Gx;
  wire   [31:0] Gy;
  tri   [7:0] OutData;
  tri   [31:0] fGy;
  tri   [31:0] fGx;
  tri   [1:0] dx;
  tri   [1:0] dy;
  tri   \regZ[0][7] ;
  tri   \regZ[0][6] ;
  tri   \regZ[0][5] ;
  tri   \regZ[0][4] ;
  tri   \regZ[0][3] ;
  tri   \regZ[0][2] ;
  tri   \regZ[0][1] ;
  tri   \regZ[0][0] ;
  tri   \regZ[1][7] ;
  tri   \regZ[1][6] ;
  tri   \regZ[1][5] ;
  tri   \regZ[1][4] ;
  tri   \regZ[1][3] ;
  tri   \regZ[1][2] ;
  tri   \regZ[1][1] ;
  tri   \regZ[1][0] ;
  tri   \regZ[2][7] ;
  tri   \regZ[2][6] ;
  tri   \regZ[2][5] ;
  tri   \regZ[2][4] ;
  tri   \regZ[2][3] ;
  tri   \regZ[2][2] ;
  tri   \regZ[2][1] ;
  tri   \regZ[2][0] ;
  tri   \regZ[3][7] ;
  tri   \regZ[3][6] ;
  tri   \regZ[3][5] ;
  tri   \regZ[3][4] ;
  tri   \regZ[3][3] ;
  tri   \regZ[3][2] ;
  tri   \regZ[3][1] ;
  tri   \regZ[3][0] ;
  tri   \regZ[4][7] ;
  tri   \regZ[4][6] ;
  tri   \regZ[4][5] ;
  tri   \regZ[4][4] ;
  tri   \regZ[4][3] ;
  tri   \regZ[4][2] ;
  tri   \regZ[4][1] ;
  tri   \regZ[4][0] ;
  tri   \regZ[5][7] ;
  tri   \regZ[5][6] ;
  tri   \regZ[5][5] ;
  tri   \regZ[5][4] ;
  tri   \regZ[5][3] ;
  tri   \regZ[5][2] ;
  tri   \regZ[5][1] ;
  tri   \regZ[5][0] ;
  tri   \regZ[6][7] ;
  tri   \regZ[6][6] ;
  tri   \regZ[6][5] ;
  tri   \regZ[6][4] ;
  tri   \regZ[6][3] ;
  tri   \regZ[6][2] ;
  tri   \regZ[6][1] ;
  tri   \regZ[6][0] ;
  tri   \regZ[7][7] ;
  tri   \regZ[7][6] ;
  tri   \regZ[7][5] ;
  tri   \regZ[7][4] ;
  tri   \regZ[7][3] ;
  tri   \regZ[7][2] ;
  tri   \regZ[7][1] ;
  tri   \regZ[7][0] ;
  tri   \regZ[8][7] ;
  tri   \regZ[8][6] ;
  tri   \regZ[8][5] ;
  tri   \regZ[8][4] ;
  tri   \regZ[8][3] ;
  tri   \regZ[8][2] ;
  tri   \regZ[8][1] ;
  tri   \regZ[8][0] ;
  tri   \regZ[9][7] ;
  tri   \regZ[9][6] ;
  tri   \regZ[9][5] ;
  tri   \regZ[9][4] ;
  tri   \regZ[9][3] ;
  tri   \regZ[9][2] ;
  tri   \regZ[9][1] ;
  tri   \regZ[9][0] ;
  tri   \regZ[10][7] ;
  tri   \regZ[10][6] ;
  tri   \regZ[10][5] ;
  tri   \regZ[10][4] ;
  tri   \regZ[10][3] ;
  tri   \regZ[10][2] ;
  tri   \regZ[10][1] ;
  tri   \regZ[10][0] ;
  tri   \regZ[11][7] ;
  tri   \regZ[11][6] ;
  tri   \regZ[11][5] ;
  tri   \regZ[11][4] ;
  tri   \regZ[11][3] ;
  tri   \regZ[11][2] ;
  tri   \regZ[11][1] ;
  tri   \regZ[11][0] ;
  tri   \regZ[12][7] ;
  tri   \regZ[12][6] ;
  tri   \regZ[12][5] ;
  tri   \regZ[12][4] ;
  tri   \regZ[12][3] ;
  tri   \regZ[12][2] ;
  tri   \regZ[12][1] ;
  tri   \regZ[12][0] ;
  tri   \regZ[13][7] ;
  tri   \regZ[13][6] ;
  tri   \regZ[13][5] ;
  tri   \regZ[13][4] ;
  tri   \regZ[13][3] ;
  tri   \regZ[13][2] ;
  tri   \regZ[13][1] ;
  tri   \regZ[13][0] ;
  tri   \regZ[14][7] ;
  tri   \regZ[14][6] ;
  tri   \regZ[14][5] ;
  tri   \regZ[14][4] ;
  tri   \regZ[14][3] ;
  tri   \regZ[14][2] ;
  tri   \regZ[14][1] ;
  tri   \regZ[14][0] ;
  tri   \regZ[15][7] ;
  tri   \regZ[15][6] ;
  tri   \regZ[15][5] ;
  tri   \regZ[15][4] ;
  tri   \regZ[15][3] ;
  tri   \regZ[15][2] ;
  tri   \regZ[15][1] ;
  tri   \regZ[15][0] ;
  tri   \regZ[16][7] ;
  tri   \regZ[16][6] ;
  tri   \regZ[16][5] ;
  tri   \regZ[16][4] ;
  tri   \regZ[16][3] ;
  tri   \regZ[16][2] ;
  tri   \regZ[16][1] ;
  tri   \regZ[16][0] ;
  tri   \regZ[17][7] ;
  tri   \regZ[17][6] ;
  tri   \regZ[17][5] ;
  tri   \regZ[17][4] ;
  tri   \regZ[17][3] ;
  tri   \regZ[17][2] ;
  tri   \regZ[17][1] ;
  tri   \regZ[17][0] ;
  tri   \regZ[18][7] ;
  tri   \regZ[18][6] ;
  tri   \regZ[18][5] ;
  tri   \regZ[18][4] ;
  tri   \regZ[18][3] ;
  tri   \regZ[18][2] ;
  tri   \regZ[18][1] ;
  tri   \regZ[18][0] ;
  tri   \regZ[19][7] ;
  tri   \regZ[19][6] ;
  tri   \regZ[19][5] ;
  tri   \regZ[19][4] ;
  tri   \regZ[19][3] ;
  tri   \regZ[19][2] ;
  tri   \regZ[19][1] ;
  tri   \regZ[19][0] ;
  tri   \regZ[20][7] ;
  tri   \regZ[20][6] ;
  tri   \regZ[20][5] ;
  tri   \regZ[20][4] ;
  tri   \regZ[20][3] ;
  tri   \regZ[20][2] ;
  tri   \regZ[20][1] ;
  tri   \regZ[20][0] ;
  tri   \regZ[21][7] ;
  tri   \regZ[21][6] ;
  tri   \regZ[21][5] ;
  tri   \regZ[21][4] ;
  tri   \regZ[21][3] ;
  tri   \regZ[21][2] ;
  tri   \regZ[21][1] ;
  tri   \regZ[21][0] ;
  tri   \regZ[22][7] ;
  tri   \regZ[22][6] ;
  tri   \regZ[22][5] ;
  tri   \regZ[22][4] ;
  tri   \regZ[22][3] ;
  tri   \regZ[22][2] ;
  tri   \regZ[22][1] ;
  tri   \regZ[22][0] ;
  tri   \regZ[23][7] ;
  tri   \regZ[23][6] ;
  tri   \regZ[23][5] ;
  tri   \regZ[23][4] ;
  tri   \regZ[23][3] ;
  tri   \regZ[23][2] ;
  tri   \regZ[23][1] ;
  tri   \regZ[23][0] ;
  tri   \regZ[24][7] ;
  tri   \regZ[24][6] ;
  tri   \regZ[24][5] ;
  tri   \regZ[24][4] ;
  tri   \regZ[24][3] ;
  tri   \regZ[24][2] ;
  tri   \regZ[24][1] ;
  tri   \regZ[24][0] ;
  tri   [7:0] Out_gradient;
  tri   [7:0] Out_direction;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80;

  DFFPOSX1 \OutData_tri_enable_reg[7]  ( .D(n5443), .CLK(clk), .Q(N4469) );
  DFFPOSX1 \OutData_tri_enable_reg[6]  ( .D(n5442), .CLK(clk), .Q(N4472) );
  DFFPOSX1 \OutData_tri_enable_reg[5]  ( .D(n5441), .CLK(clk), .Q(N4475) );
  DFFPOSX1 \OutData_tri_enable_reg[4]  ( .D(n5440), .CLK(clk), .Q(N4478) );
  DFFPOSX1 \OutData_tri_enable_reg[3]  ( .D(n5439), .CLK(clk), .Q(N4481) );
  DFFPOSX1 \OutData_tri_enable_reg[2]  ( .D(n5438), .CLK(clk), .Q(N4484) );
  DFFPOSX1 \OutData_tri_enable_reg[1]  ( .D(n5437), .CLK(clk), .Q(N4487) );
  DFFPOSX1 \OutData_tri_enable_reg[0]  ( .D(n5436), .CLK(clk), .Q(N4490) );
  DFFSR \IntSignal_reg[0]  ( .D(n5435), .CLK(clk), .R(rst_b), .S(1'b1), .Q(
        IntSignal[0]) );
  DFFSR \IntSignal_reg[1]  ( .D(n5434), .CLK(clk), .R(rst_b), .S(1'b1), .Q(
        IntSignal[1]) );
  DFFPOSX1 \fGx_tri_enable_reg[0]  ( .D(n5433), .CLK(clk), .Q(N4394) );
  DFFPOSX1 \fGx_tri_enable_reg[1]  ( .D(n5432), .CLK(clk), .Q(N4391) );
  DFFPOSX1 \fGx_tri_enable_reg[2]  ( .D(n5431), .CLK(clk), .Q(N4388) );
  DFFPOSX1 \fGx_tri_enable_reg[3]  ( .D(n5430), .CLK(clk), .Q(N4385) );
  DFFPOSX1 \fGx_tri_enable_reg[4]  ( .D(n5429), .CLK(clk), .Q(N4382) );
  DFFPOSX1 \fGx_tri_enable_reg[5]  ( .D(n5428), .CLK(clk), .Q(N4379) );
  DFFPOSX1 \fGx_tri_enable_reg[6]  ( .D(n5427), .CLK(clk), .Q(N4376) );
  DFFPOSX1 \fGx_tri_enable_reg[7]  ( .D(n5426), .CLK(clk), .Q(N4373) );
  DFFPOSX1 \fGy_tri_enable_reg[0]  ( .D(n5425), .CLK(clk), .Q(N4466) );
  DFFPOSX1 \fGy_tri_enable_reg[1]  ( .D(n5424), .CLK(clk), .Q(N4463) );
  DFFPOSX1 \fGy_tri_enable_reg[2]  ( .D(n5423), .CLK(clk), .Q(N4460) );
  DFFPOSX1 \fGy_tri_enable_reg[3]  ( .D(n5422), .CLK(clk), .Q(N4457) );
  DFFPOSX1 \fGy_tri_enable_reg[4]  ( .D(n5421), .CLK(clk), .Q(N4454) );
  DFFPOSX1 \fGy_tri_enable_reg[5]  ( .D(n5420), .CLK(clk), .Q(N4451) );
  DFFPOSX1 \fGy_tri_enable_reg[6]  ( .D(n5419), .CLK(clk), .Q(N4448) );
  DFFPOSX1 \fGy_tri_enable_reg[7]  ( .D(n5418), .CLK(clk), .Q(N4445) );
  DFFPOSX1 \dx_tri_enable_reg[0]  ( .D(n5417), .CLK(clk), .Q(N4502) );
  DFFPOSX1 \regX_reg[15][0]  ( .D(n5344), .CLK(clk), .Q(\regX[15][0] ) );
  DFFPOSX1 \regX_reg[15][1]  ( .D(n5343), .CLK(clk), .Q(\regX[15][1] ) );
  DFFPOSX1 \regX_reg[15][2]  ( .D(n5342), .CLK(clk), .Q(\regX[15][2] ) );
  DFFPOSX1 \regX_reg[15][3]  ( .D(n5341), .CLK(clk), .Q(\regX[15][3] ) );
  DFFPOSX1 \regX_reg[15][4]  ( .D(n5340), .CLK(clk), .Q(\regX[15][4] ) );
  DFFPOSX1 \regX_reg[15][5]  ( .D(n5339), .CLK(clk), .Q(\regX[15][5] ) );
  DFFPOSX1 \regX_reg[15][6]  ( .D(n5338), .CLK(clk), .Q(\regX[15][6] ) );
  DFFPOSX1 \regX_reg[15][7]  ( .D(n5337), .CLK(clk), .Q(\regX[15][7] ) );
  DFFPOSX1 \regX_reg[1][0]  ( .D(n5232), .CLK(clk), .Q(\regX[1][0] ) );
  DFFPOSX1 \regX_reg[1][1]  ( .D(n5231), .CLK(clk), .Q(\regX[1][1] ) );
  DFFPOSX1 \regX_reg[1][2]  ( .D(n5230), .CLK(clk), .Q(\regX[1][2] ) );
  DFFPOSX1 \regX_reg[1][3]  ( .D(n5229), .CLK(clk), .Q(\regX[1][3] ) );
  DFFPOSX1 \regX_reg[1][4]  ( .D(n5228), .CLK(clk), .Q(\regX[1][4] ) );
  DFFPOSX1 \regX_reg[1][5]  ( .D(n5227), .CLK(clk), .Q(\regX[1][5] ) );
  DFFPOSX1 \regX_reg[1][6]  ( .D(n5226), .CLK(clk), .Q(\regX[1][6] ) );
  DFFPOSX1 \regX_reg[1][7]  ( .D(n5225), .CLK(clk), .Q(\regX[1][7] ) );
  DFFPOSX1 \regX_reg[24][0]  ( .D(n5416), .CLK(clk), .Q(\regX[24][0] ) );
  DFFPOSX1 \regX_reg[24][1]  ( .D(n5415), .CLK(clk), .Q(\regX[24][1] ) );
  DFFPOSX1 \regX_reg[24][2]  ( .D(n5414), .CLK(clk), .Q(\regX[24][2] ) );
  DFFPOSX1 \regX_reg[24][3]  ( .D(n5413), .CLK(clk), .Q(\regX[24][3] ) );
  DFFPOSX1 \regX_reg[24][4]  ( .D(n5412), .CLK(clk), .Q(\regX[24][4] ) );
  DFFPOSX1 \regX_reg[24][5]  ( .D(n5411), .CLK(clk), .Q(\regX[24][5] ) );
  DFFPOSX1 \regX_reg[24][6]  ( .D(n5410), .CLK(clk), .Q(\regX[24][6] ) );
  DFFPOSX1 \regX_reg[24][7]  ( .D(n5409), .CLK(clk), .Q(\regX[24][7] ) );
  DFFPOSX1 \regX_reg[16][0]  ( .D(n5352), .CLK(clk), .Q(\regX[16][0] ) );
  DFFPOSX1 \regX_reg[16][1]  ( .D(n5351), .CLK(clk), .Q(\regX[16][1] ) );
  DFFPOSX1 \regX_reg[16][2]  ( .D(n5350), .CLK(clk), .Q(\regX[16][2] ) );
  DFFPOSX1 \regX_reg[16][3]  ( .D(n5349), .CLK(clk), .Q(\regX[16][3] ) );
  DFFPOSX1 \regX_reg[16][4]  ( .D(n5348), .CLK(clk), .Q(\regX[16][4] ) );
  DFFPOSX1 \regX_reg[16][5]  ( .D(n5347), .CLK(clk), .Q(\regX[16][5] ) );
  DFFPOSX1 \regX_reg[16][6]  ( .D(n5346), .CLK(clk), .Q(\regX[16][6] ) );
  DFFPOSX1 \regX_reg[16][7]  ( .D(n5345), .CLK(clk), .Q(\regX[16][7] ) );
  DFFPOSX1 \regX_reg[17][0]  ( .D(n5360), .CLK(clk), .Q(\regX[17][0] ) );
  DFFPOSX1 \regX_reg[17][1]  ( .D(n5359), .CLK(clk), .Q(\regX[17][1] ) );
  DFFPOSX1 \regX_reg[17][2]  ( .D(n5358), .CLK(clk), .Q(\regX[17][2] ) );
  DFFPOSX1 \regX_reg[17][3]  ( .D(n5357), .CLK(clk), .Q(\regX[17][3] ) );
  DFFPOSX1 \regX_reg[17][4]  ( .D(n5356), .CLK(clk), .Q(\regX[17][4] ) );
  DFFPOSX1 \regX_reg[17][5]  ( .D(n5355), .CLK(clk), .Q(\regX[17][5] ) );
  DFFPOSX1 \regX_reg[17][6]  ( .D(n5354), .CLK(clk), .Q(\regX[17][6] ) );
  DFFPOSX1 \regX_reg[17][7]  ( .D(n5353), .CLK(clk), .Q(\regX[17][7] ) );
  DFFPOSX1 \regX_reg[18][0]  ( .D(n5368), .CLK(clk), .Q(\regX[18][0] ) );
  DFFPOSX1 \regX_reg[18][1]  ( .D(n5367), .CLK(clk), .Q(\regX[18][1] ) );
  DFFPOSX1 \regX_reg[18][2]  ( .D(n5366), .CLK(clk), .Q(\regX[18][2] ) );
  DFFPOSX1 \regX_reg[18][3]  ( .D(n5365), .CLK(clk), .Q(\regX[18][3] ) );
  DFFPOSX1 \regX_reg[18][4]  ( .D(n5364), .CLK(clk), .Q(\regX[18][4] ) );
  DFFPOSX1 \regX_reg[18][5]  ( .D(n5363), .CLK(clk), .Q(\regX[18][5] ) );
  DFFPOSX1 \regX_reg[18][6]  ( .D(n5362), .CLK(clk), .Q(\regX[18][6] ) );
  DFFPOSX1 \regX_reg[18][7]  ( .D(n5361), .CLK(clk), .Q(\regX[18][7] ) );
  DFFPOSX1 \regX_reg[20][0]  ( .D(n5384), .CLK(clk), .Q(\regX[20][0] ) );
  DFFPOSX1 \regX_reg[20][1]  ( .D(n5383), .CLK(clk), .Q(\regX[20][1] ) );
  DFFPOSX1 \regX_reg[20][2]  ( .D(n5382), .CLK(clk), .Q(\regX[20][2] ) );
  DFFPOSX1 \regX_reg[20][3]  ( .D(n5381), .CLK(clk), .Q(\regX[20][3] ) );
  DFFPOSX1 \regX_reg[20][4]  ( .D(n5380), .CLK(clk), .Q(\regX[20][4] ) );
  DFFPOSX1 \regX_reg[20][5]  ( .D(n5379), .CLK(clk), .Q(\regX[20][5] ) );
  DFFPOSX1 \regX_reg[20][6]  ( .D(n5378), .CLK(clk), .Q(\regX[20][6] ) );
  DFFPOSX1 \regX_reg[20][7]  ( .D(n5377), .CLK(clk), .Q(\regX[20][7] ) );
  DFFPOSX1 \regX_reg[22][0]  ( .D(n5400), .CLK(clk), .Q(\regX[22][0] ) );
  DFFPOSX1 \regX_reg[22][1]  ( .D(n5399), .CLK(clk), .Q(\regX[22][1] ) );
  DFFPOSX1 \regX_reg[22][2]  ( .D(n5398), .CLK(clk), .Q(\regX[22][2] ) );
  DFFPOSX1 \regX_reg[22][3]  ( .D(n5397), .CLK(clk), .Q(\regX[22][3] ) );
  DFFPOSX1 \regX_reg[22][4]  ( .D(n5396), .CLK(clk), .Q(\regX[22][4] ) );
  DFFPOSX1 \regX_reg[22][5]  ( .D(n5395), .CLK(clk), .Q(\regX[22][5] ) );
  DFFPOSX1 \regX_reg[22][6]  ( .D(n5394), .CLK(clk), .Q(\regX[22][6] ) );
  DFFPOSX1 \regX_reg[22][7]  ( .D(n5393), .CLK(clk), .Q(\regX[22][7] ) );
  DFFPOSX1 \regX_reg[19][0]  ( .D(n5376), .CLK(clk), .Q(\regX[19][0] ) );
  DFFPOSX1 \regX_reg[19][1]  ( .D(n5375), .CLK(clk), .Q(\regX[19][1] ) );
  DFFPOSX1 \regX_reg[19][2]  ( .D(n5374), .CLK(clk), .Q(\regX[19][2] ) );
  DFFPOSX1 \regX_reg[19][3]  ( .D(n5373), .CLK(clk), .Q(\regX[19][3] ) );
  DFFPOSX1 \regX_reg[19][4]  ( .D(n5372), .CLK(clk), .Q(\regX[19][4] ) );
  DFFPOSX1 \regX_reg[19][5]  ( .D(n5371), .CLK(clk), .Q(\regX[19][5] ) );
  DFFPOSX1 \regX_reg[19][6]  ( .D(n5370), .CLK(clk), .Q(\regX[19][6] ) );
  DFFPOSX1 \regX_reg[19][7]  ( .D(n5369), .CLK(clk), .Q(\regX[19][7] ) );
  DFFPOSX1 \regX_reg[21][0]  ( .D(n5392), .CLK(clk), .Q(\regX[21][0] ) );
  DFFPOSX1 \regX_reg[21][1]  ( .D(n5391), .CLK(clk), .Q(\regX[21][1] ) );
  DFFPOSX1 \regX_reg[21][2]  ( .D(n5390), .CLK(clk), .Q(\regX[21][2] ) );
  DFFPOSX1 \regX_reg[21][3]  ( .D(n5389), .CLK(clk), .Q(\regX[21][3] ) );
  DFFPOSX1 \regX_reg[21][4]  ( .D(n5388), .CLK(clk), .Q(\regX[21][4] ) );
  DFFPOSX1 \regX_reg[21][5]  ( .D(n5387), .CLK(clk), .Q(\regX[21][5] ) );
  DFFPOSX1 \regX_reg[21][6]  ( .D(n5386), .CLK(clk), .Q(\regX[21][6] ) );
  DFFPOSX1 \regX_reg[21][7]  ( .D(n5385), .CLK(clk), .Q(\regX[21][7] ) );
  DFFPOSX1 \regX_reg[23][0]  ( .D(n5408), .CLK(clk), .Q(\regX[23][0] ) );
  DFFPOSX1 \regX_reg[23][1]  ( .D(n5407), .CLK(clk), .Q(\regX[23][1] ) );
  DFFPOSX1 \regX_reg[23][2]  ( .D(n5406), .CLK(clk), .Q(\regX[23][2] ) );
  DFFPOSX1 \regX_reg[23][3]  ( .D(n5405), .CLK(clk), .Q(\regX[23][3] ) );
  DFFPOSX1 \regX_reg[23][4]  ( .D(n5404), .CLK(clk), .Q(\regX[23][4] ) );
  DFFPOSX1 \regX_reg[23][5]  ( .D(n5403), .CLK(clk), .Q(\regX[23][5] ) );
  DFFPOSX1 \regX_reg[23][6]  ( .D(n5402), .CLK(clk), .Q(\regX[23][6] ) );
  DFFPOSX1 \regX_reg[23][7]  ( .D(n5401), .CLK(clk), .Q(\regX[23][7] ) );
  DFFPOSX1 \regX_reg[8][0]  ( .D(n5288), .CLK(clk), .Q(\regX[8][0] ) );
  DFFPOSX1 \regX_reg[8][1]  ( .D(n5287), .CLK(clk), .Q(\regX[8][1] ) );
  DFFPOSX1 \regX_reg[8][2]  ( .D(n5286), .CLK(clk), .Q(\regX[8][2] ) );
  DFFPOSX1 \regX_reg[8][3]  ( .D(n5285), .CLK(clk), .Q(\regX[8][3] ) );
  DFFPOSX1 \regX_reg[8][4]  ( .D(n5284), .CLK(clk), .Q(\regX[8][4] ) );
  DFFPOSX1 \regX_reg[8][5]  ( .D(n5283), .CLK(clk), .Q(\regX[8][5] ) );
  DFFPOSX1 \regX_reg[8][6]  ( .D(n5282), .CLK(clk), .Q(\regX[8][6] ) );
  DFFPOSX1 \regX_reg[8][7]  ( .D(n5281), .CLK(clk), .Q(\regX[8][7] ) );
  DFFPOSX1 \regX_reg[9][0]  ( .D(n5296), .CLK(clk), .Q(\regX[9][0] ) );
  DFFPOSX1 \regX_reg[9][1]  ( .D(n5295), .CLK(clk), .Q(\regX[9][1] ) );
  DFFPOSX1 \regX_reg[9][2]  ( .D(n5294), .CLK(clk), .Q(\regX[9][2] ) );
  DFFPOSX1 \regX_reg[9][3]  ( .D(n5293), .CLK(clk), .Q(\regX[9][3] ) );
  DFFPOSX1 \regX_reg[9][4]  ( .D(n5292), .CLK(clk), .Q(\regX[9][4] ) );
  DFFPOSX1 \regX_reg[9][5]  ( .D(n5291), .CLK(clk), .Q(\regX[9][5] ) );
  DFFPOSX1 \regX_reg[9][6]  ( .D(n5290), .CLK(clk), .Q(\regX[9][6] ) );
  DFFPOSX1 \regX_reg[9][7]  ( .D(n5289), .CLK(clk), .Q(\regX[9][7] ) );
  DFFPOSX1 \regX_reg[10][0]  ( .D(n5304), .CLK(clk), .Q(N1615) );
  DFFPOSX1 \regX_reg[10][1]  ( .D(n5303), .CLK(clk), .Q(N1616) );
  DFFPOSX1 \regX_reg[10][2]  ( .D(n5302), .CLK(clk), .Q(N1617) );
  DFFPOSX1 \regX_reg[10][3]  ( .D(n5301), .CLK(clk), .Q(N1618) );
  DFFPOSX1 \regX_reg[10][4]  ( .D(n5300), .CLK(clk), .Q(N1619) );
  DFFPOSX1 \regX_reg[10][5]  ( .D(n5299), .CLK(clk), .Q(N1620) );
  DFFPOSX1 \regX_reg[10][6]  ( .D(n5298), .CLK(clk), .Q(N1621) );
  DFFPOSX1 \regX_reg[10][7]  ( .D(n5297), .CLK(clk), .Q(N1622) );
  DFFPOSX1 \regX_reg[12][0]  ( .D(n5320), .CLK(clk), .Q(N1677) );
  DFFPOSX1 \regX_reg[12][1]  ( .D(n5319), .CLK(clk), .Q(N1678) );
  DFFPOSX1 \regX_reg[12][2]  ( .D(n5318), .CLK(clk), .Q(N1679) );
  DFFPOSX1 \regX_reg[12][3]  ( .D(n5317), .CLK(clk), .Q(N1680) );
  DFFPOSX1 \regX_reg[12][4]  ( .D(n5316), .CLK(clk), .Q(N1681) );
  DFFPOSX1 \regX_reg[12][5]  ( .D(n5315), .CLK(clk), .Q(N1682) );
  DFFPOSX1 \regX_reg[12][6]  ( .D(n5314), .CLK(clk), .Q(N1683) );
  DFFPOSX1 \regX_reg[12][7]  ( .D(n5313), .CLK(clk), .Q(N1684) );
  DFFPOSX1 \regX_reg[14][0]  ( .D(n5336), .CLK(clk), .Q(N1735) );
  DFFPOSX1 \regX_reg[14][1]  ( .D(n5335), .CLK(clk), .Q(N1736) );
  DFFPOSX1 \regX_reg[14][2]  ( .D(n5334), .CLK(clk), .Q(N1737) );
  DFFPOSX1 \regX_reg[14][3]  ( .D(n5333), .CLK(clk), .Q(N1738) );
  DFFPOSX1 \regX_reg[14][4]  ( .D(n5332), .CLK(clk), .Q(N1739) );
  DFFPOSX1 \regX_reg[14][5]  ( .D(n5331), .CLK(clk), .Q(N1740) );
  DFFPOSX1 \regX_reg[14][6]  ( .D(n5330), .CLK(clk), .Q(N1741) );
  DFFPOSX1 \regX_reg[14][7]  ( .D(n5329), .CLK(clk), .Q(N1742) );
  DFFPOSX1 \regX_reg[11][0]  ( .D(n5312), .CLK(clk), .Q(\regX[11][0] ) );
  DFFPOSX1 \regX_reg[11][1]  ( .D(n5311), .CLK(clk), .Q(\regX[11][1] ) );
  DFFPOSX1 \regX_reg[11][2]  ( .D(n5310), .CLK(clk), .Q(\regX[11][2] ) );
  DFFPOSX1 \regX_reg[11][3]  ( .D(n5309), .CLK(clk), .Q(\regX[11][3] ) );
  DFFPOSX1 \regX_reg[11][4]  ( .D(n5308), .CLK(clk), .Q(\regX[11][4] ) );
  DFFPOSX1 \regX_reg[11][5]  ( .D(n5307), .CLK(clk), .Q(\regX[11][5] ) );
  DFFPOSX1 \regX_reg[11][6]  ( .D(n5306), .CLK(clk), .Q(\regX[11][6] ) );
  DFFPOSX1 \regX_reg[11][7]  ( .D(n5305), .CLK(clk), .Q(\regX[11][7] ) );
  DFFPOSX1 \regX_reg[2][0]  ( .D(n5240), .CLK(clk), .Q(N1375) );
  DFFPOSX1 \regX_reg[2][1]  ( .D(n5239), .CLK(clk), .Q(N1376) );
  DFFPOSX1 \regX_reg[2][2]  ( .D(n5238), .CLK(clk), .Q(N1377) );
  DFFPOSX1 \regX_reg[2][3]  ( .D(n5237), .CLK(clk), .Q(N1378) );
  DFFPOSX1 \regX_reg[2][4]  ( .D(n5236), .CLK(clk), .Q(N1379) );
  DFFPOSX1 \regX_reg[2][5]  ( .D(n5235), .CLK(clk), .Q(N1380) );
  DFFPOSX1 \regX_reg[2][6]  ( .D(n5234), .CLK(clk), .Q(N1381) );
  DFFPOSX1 \regX_reg[2][7]  ( .D(n5233), .CLK(clk), .Q(N1382) );
  DFFPOSX1 \regX_reg[4][0]  ( .D(n5256), .CLK(clk), .Q(N1433) );
  DFFPOSX1 \regX_reg[4][1]  ( .D(n5255), .CLK(clk), .Q(N1434) );
  DFFPOSX1 \regX_reg[4][2]  ( .D(n5254), .CLK(clk), .Q(N1435) );
  DFFPOSX1 \regX_reg[4][3]  ( .D(n5253), .CLK(clk), .Q(N1436) );
  DFFPOSX1 \regX_reg[4][4]  ( .D(n5252), .CLK(clk), .Q(N1437) );
  DFFPOSX1 \regX_reg[4][5]  ( .D(n5251), .CLK(clk), .Q(N1438) );
  DFFPOSX1 \regX_reg[4][6]  ( .D(n5250), .CLK(clk), .Q(N1439) );
  DFFPOSX1 \regX_reg[4][7]  ( .D(n5249), .CLK(clk), .Q(N1440) );
  DFFPOSX1 \regX_reg[3][0]  ( .D(n5248), .CLK(clk), .Q(\regX[3][0] ) );
  DFFPOSX1 \regX_reg[3][1]  ( .D(n5247), .CLK(clk), .Q(\regX[3][1] ) );
  DFFPOSX1 \regX_reg[3][2]  ( .D(n5246), .CLK(clk), .Q(\regX[3][2] ) );
  DFFPOSX1 \regX_reg[3][3]  ( .D(n5245), .CLK(clk), .Q(\regX[3][3] ) );
  DFFPOSX1 \regX_reg[3][4]  ( .D(n5244), .CLK(clk), .Q(\regX[3][4] ) );
  DFFPOSX1 \regX_reg[3][5]  ( .D(n5243), .CLK(clk), .Q(\regX[3][5] ) );
  DFFPOSX1 \regX_reg[3][6]  ( .D(n5242), .CLK(clk), .Q(\regX[3][6] ) );
  DFFPOSX1 \regX_reg[3][7]  ( .D(n5241), .CLK(clk), .Q(\regX[3][7] ) );
  DFFPOSX1 \regX_reg[5][0]  ( .D(n5264), .CLK(clk), .Q(\regX[5][0] ) );
  DFFPOSX1 \regX_reg[5][1]  ( .D(n5263), .CLK(clk), .Q(\regX[5][1] ) );
  DFFPOSX1 \regX_reg[5][2]  ( .D(n5262), .CLK(clk), .Q(\regX[5][2] ) );
  DFFPOSX1 \regX_reg[5][3]  ( .D(n5261), .CLK(clk), .Q(\regX[5][3] ) );
  DFFPOSX1 \regX_reg[5][4]  ( .D(n5260), .CLK(clk), .Q(\regX[5][4] ) );
  DFFPOSX1 \regX_reg[5][5]  ( .D(n5259), .CLK(clk), .Q(\regX[5][5] ) );
  DFFPOSX1 \regX_reg[5][6]  ( .D(n5258), .CLK(clk), .Q(\regX[5][6] ) );
  DFFPOSX1 \regX_reg[5][7]  ( .D(n5257), .CLK(clk), .Q(\regX[5][7] ) );
  DFFPOSX1 \regX_reg[7][0]  ( .D(n5280), .CLK(clk), .Q(\regX[7][0] ) );
  DFFPOSX1 \regX_reg[7][1]  ( .D(n5279), .CLK(clk), .Q(\regX[7][1] ) );
  DFFPOSX1 \regX_reg[7][2]  ( .D(n5278), .CLK(clk), .Q(\regX[7][2] ) );
  DFFPOSX1 \regX_reg[7][3]  ( .D(n5277), .CLK(clk), .Q(\regX[7][3] ) );
  DFFPOSX1 \regX_reg[7][4]  ( .D(n5276), .CLK(clk), .Q(\regX[7][4] ) );
  DFFPOSX1 \regX_reg[7][5]  ( .D(n5275), .CLK(clk), .Q(\regX[7][5] ) );
  DFFPOSX1 \regX_reg[7][6]  ( .D(n5274), .CLK(clk), .Q(\regX[7][6] ) );
  DFFPOSX1 \regX_reg[7][7]  ( .D(n5273), .CLK(clk), .Q(\regX[7][7] ) );
  DFFPOSX1 \regX_reg[13][7]  ( .D(n5328), .CLK(clk), .Q(\regX[13][7] ) );
  DFFPOSX1 \regX_reg[13][0]  ( .D(n5327), .CLK(clk), .Q(\regX[13][0] ) );
  DFFPOSX1 \regX_reg[13][1]  ( .D(n5326), .CLK(clk), .Q(\regX[13][1] ) );
  DFFPOSX1 \regX_reg[13][2]  ( .D(n5325), .CLK(clk), .Q(\regX[13][2] ) );
  DFFPOSX1 \regX_reg[13][3]  ( .D(n5324), .CLK(clk), .Q(\regX[13][3] ) );
  DFFPOSX1 \regX_reg[13][4]  ( .D(n5323), .CLK(clk), .Q(\regX[13][4] ) );
  DFFPOSX1 \regX_reg[13][5]  ( .D(n5322), .CLK(clk), .Q(\regX[13][5] ) );
  DFFPOSX1 \regX_reg[13][6]  ( .D(n5321), .CLK(clk), .Q(\regX[13][6] ) );
  DFFPOSX1 \regY_reg[6][0]  ( .D(n3682), .CLK(clk), .Q(\regY[6][0] ) );
  DFFPOSX1 \regY_reg[6][1]  ( .D(n3683), .CLK(clk), .Q(\regY[6][1] ) );
  DFFPOSX1 \regY_reg[6][2]  ( .D(n3684), .CLK(clk), .Q(\regY[6][2] ) );
  DFFPOSX1 \regY_reg[6][3]  ( .D(n3685), .CLK(clk), .Q(\regY[6][3] ) );
  DFFPOSX1 \regY_reg[6][4]  ( .D(n3686), .CLK(clk), .Q(\regY[6][4] ) );
  DFFPOSX1 \regY_reg[6][5]  ( .D(n3687), .CLK(clk), .Q(\regY[6][5] ) );
  DFFPOSX1 \regY_reg[6][6]  ( .D(n7200), .CLK(clk), .Q(\regY[6][6] ) );
  DFFPOSX1 \regY_reg[6][7]  ( .D(n3688), .CLK(clk), .Q(\regY[6][7] ) );
  DFFPOSX1 \dy_reg[1]  ( .D(n4679), .CLK(clk), .Q(dy[1]) );
  DFFPOSX1 \dx_reg[1]  ( .D(n4677), .CLK(clk), .Q(dx[1]) );
  DFFPOSX1 \dx_reg[0]  ( .D(n4678), .CLK(clk), .Q(N4501) );
  DFFPOSX1 \dy_reg[0]  ( .D(n4680), .CLK(clk), .Q(N4495) );
  DFFPOSX1 \dy_tri_enable_reg[0]  ( .D(n4681), .CLK(clk), .Q(N4496) );
  DFFPOSX1 \regX_reg[6][0]  ( .D(n5272), .CLK(clk), .Q(\regX[6][0] ) );
  DFFPOSX1 \regX_reg[6][1]  ( .D(n5271), .CLK(clk), .Q(\regX[6][1] ) );
  DFFPOSX1 \regX_reg[6][2]  ( .D(n5270), .CLK(clk), .Q(\regX[6][2] ) );
  DFFPOSX1 \regX_reg[6][3]  ( .D(n5269), .CLK(clk), .Q(\regX[6][3] ) );
  DFFPOSX1 \regX_reg[6][4]  ( .D(n5268), .CLK(clk), .Q(\regX[6][4] ) );
  DFFPOSX1 \regX_reg[6][5]  ( .D(n5267), .CLK(clk), .Q(\regX[6][5] ) );
  DFFPOSX1 \regX_reg[6][6]  ( .D(n5266), .CLK(clk), .Q(\regX[6][6] ) );
  DFFPOSX1 \regX_reg[6][7]  ( .D(n5265), .CLK(clk), .Q(\regX[6][7] ) );
  DFFPOSX1 \regX_reg[0][2]  ( .D(n5224), .CLK(clk), .Q(\regX[0][2] ) );
  DFFPOSX1 \regX_reg[0][3]  ( .D(n5223), .CLK(clk), .Q(\regX[0][3] ) );
  DFFPOSX1 \regX_reg[0][4]  ( .D(n5222), .CLK(clk), .Q(\regX[0][4] ) );
  DFFPOSX1 \regX_reg[0][5]  ( .D(n5221), .CLK(clk), .Q(\regX[0][5] ) );
  DFFPOSX1 \regX_reg[0][6]  ( .D(n5220), .CLK(clk), .Q(\regX[0][6] ) );
  DFFPOSX1 \regX_reg[0][7]  ( .D(n5219), .CLK(clk), .Q(\regX[0][7] ) );
  DFFPOSX1 \regX_reg[0][0]  ( .D(n5218), .CLK(clk), .Q(\regX[0][0] ) );
  DFFPOSX1 \regX_reg[0][1]  ( .D(n5217), .CLK(clk), .Q(\regX[0][1] ) );
  DFFPOSX1 \Gy_reg[0]  ( .D(n5216), .CLK(clk), .Q(Gy[0]) );
  DFFPOSX1 \Gy_reg[1]  ( .D(n5215), .CLK(clk), .Q(Gy[1]) );
  DFFPOSX1 \Gy_reg[2]  ( .D(n5214), .CLK(clk), .Q(Gy[2]) );
  DFFPOSX1 \Gy_reg[3]  ( .D(n5213), .CLK(clk), .Q(Gy[3]) );
  DFFPOSX1 \Gy_reg[4]  ( .D(n5212), .CLK(clk), .Q(Gy[4]) );
  DFFPOSX1 \Gy_reg[5]  ( .D(n5211), .CLK(clk), .Q(Gy[5]) );
  DFFPOSX1 \Gy_reg[6]  ( .D(n5210), .CLK(clk), .Q(Gy[6]) );
  DFFPOSX1 \Gy_reg[7]  ( .D(n5209), .CLK(clk), .Q(Gy[7]) );
  DFFPOSX1 \Gy_reg[8]  ( .D(n5208), .CLK(clk), .Q(Gy[8]) );
  DFFPOSX1 \Gy_reg[9]  ( .D(n5207), .CLK(clk), .Q(Gy[9]) );
  DFFPOSX1 \Gy_reg[10]  ( .D(n5206), .CLK(clk), .Q(Gy[10]) );
  DFFPOSX1 \Gy_reg[11]  ( .D(n5205), .CLK(clk), .Q(Gy[11]) );
  DFFPOSX1 \Gy_reg[12]  ( .D(n5204), .CLK(clk), .Q(Gy[12]) );
  DFFPOSX1 \Gy_reg[13]  ( .D(n5203), .CLK(clk), .Q(Gy[13]) );
  DFFPOSX1 \Gy_reg[14]  ( .D(n5202), .CLK(clk), .Q(Gy[14]) );
  DFFPOSX1 \Gy_reg[15]  ( .D(n5201), .CLK(clk), .Q(Gy[15]) );
  DFFPOSX1 \Gy_reg[16]  ( .D(n5200), .CLK(clk), .Q(Gy[16]) );
  DFFPOSX1 \Gy_reg[17]  ( .D(n5199), .CLK(clk), .Q(Gy[17]) );
  DFFPOSX1 \Gy_reg[18]  ( .D(n5198), .CLK(clk), .Q(Gy[18]) );
  DFFPOSX1 \Gy_reg[19]  ( .D(n5197), .CLK(clk), .Q(Gy[19]) );
  DFFPOSX1 \Gy_reg[20]  ( .D(n5196), .CLK(clk), .Q(Gy[20]) );
  DFFPOSX1 \Gy_reg[21]  ( .D(n5195), .CLK(clk), .Q(Gy[21]) );
  DFFPOSX1 \Gy_reg[22]  ( .D(n5194), .CLK(clk), .Q(Gy[22]) );
  DFFPOSX1 \Gy_reg[23]  ( .D(n5193), .CLK(clk), .Q(Gy[23]) );
  DFFPOSX1 \Gy_reg[24]  ( .D(n5192), .CLK(clk), .Q(Gy[24]) );
  DFFPOSX1 \Gy_reg[25]  ( .D(n5191), .CLK(clk), .Q(Gy[25]) );
  DFFPOSX1 \Gy_reg[26]  ( .D(n5190), .CLK(clk), .Q(Gy[26]) );
  DFFPOSX1 \Gy_reg[27]  ( .D(n5189), .CLK(clk), .Q(Gy[27]) );
  DFFPOSX1 \Gy_reg[28]  ( .D(n5188), .CLK(clk), .Q(Gy[28]) );
  DFFPOSX1 \Gy_reg[29]  ( .D(n5187), .CLK(clk), .Q(Gy[29]) );
  DFFPOSX1 \Gy_reg[30]  ( .D(n5186), .CLK(clk), .Q(Gy[30]) );
  DFFPOSX1 \Gy_reg[31]  ( .D(n5185), .CLK(clk), .Q(Gy[31]) );
  DFFPOSX1 \fGx_reg[0]  ( .D(n5152), .CLK(clk), .Q(N4393) );
  DFFPOSX1 \fGy_reg[0]  ( .D(n5120), .CLK(clk), .Q(N4465) );
  DFFPOSX1 \fGy_reg[1]  ( .D(n5119), .CLK(clk), .Q(N4462) );
  DFFPOSX1 \fGy_reg[2]  ( .D(n5118), .CLK(clk), .Q(N4459) );
  DFFPOSX1 \fGy_reg[3]  ( .D(n5117), .CLK(clk), .Q(N4456) );
  DFFPOSX1 \fGy_reg[4]  ( .D(n5116), .CLK(clk), .Q(N4453) );
  DFFPOSX1 \fGy_reg[5]  ( .D(n5115), .CLK(clk), .Q(N4450) );
  DFFPOSX1 \fGy_reg[6]  ( .D(n5114), .CLK(clk), .Q(N4447) );
  DFFPOSX1 \fGy_reg[7]  ( .D(n5113), .CLK(clk), .Q(N4444) );
  DFFPOSX1 \fGy_reg[8]  ( .D(n5112), .CLK(clk), .Q(fGy[8]) );
  DFFPOSX1 \fGy_reg[9]  ( .D(n5111), .CLK(clk), .Q(fGy[9]) );
  DFFPOSX1 \fGy_reg[10]  ( .D(n5110), .CLK(clk), .Q(fGy[10]) );
  DFFPOSX1 \fGy_reg[11]  ( .D(n5109), .CLK(clk), .Q(fGy[11]) );
  DFFPOSX1 \fGy_reg[12]  ( .D(n5108), .CLK(clk), .Q(fGy[12]) );
  DFFPOSX1 \fGy_reg[13]  ( .D(n5107), .CLK(clk), .Q(fGy[13]) );
  DFFPOSX1 \fGy_reg[14]  ( .D(n5106), .CLK(clk), .Q(fGy[14]) );
  DFFPOSX1 \fGy_reg[15]  ( .D(n5105), .CLK(clk), .Q(fGy[15]) );
  DFFPOSX1 \fGy_reg[16]  ( .D(n5104), .CLK(clk), .Q(fGy[16]) );
  DFFPOSX1 \fGy_reg[17]  ( .D(n5103), .CLK(clk), .Q(fGy[17]) );
  DFFPOSX1 \fGy_reg[18]  ( .D(n5102), .CLK(clk), .Q(fGy[18]) );
  DFFPOSX1 \fGy_reg[19]  ( .D(n5101), .CLK(clk), .Q(fGy[19]) );
  DFFPOSX1 \fGy_reg[20]  ( .D(n5100), .CLK(clk), .Q(fGy[20]) );
  DFFPOSX1 \fGy_reg[21]  ( .D(n5099), .CLK(clk), .Q(fGy[21]) );
  DFFPOSX1 \fGy_reg[22]  ( .D(n5098), .CLK(clk), .Q(fGy[22]) );
  DFFPOSX1 \fGy_reg[23]  ( .D(n5097), .CLK(clk), .Q(fGy[23]) );
  DFFPOSX1 \fGy_reg[24]  ( .D(n5096), .CLK(clk), .Q(fGy[24]) );
  DFFPOSX1 \fGy_reg[25]  ( .D(n5095), .CLK(clk), .Q(fGy[25]) );
  DFFPOSX1 \fGy_reg[26]  ( .D(n5094), .CLK(clk), .Q(fGy[26]) );
  DFFPOSX1 \fGy_reg[27]  ( .D(n5093), .CLK(clk), .Q(fGy[27]) );
  DFFPOSX1 \fGy_reg[28]  ( .D(n5092), .CLK(clk), .Q(fGy[28]) );
  DFFPOSX1 \fGy_reg[29]  ( .D(n5091), .CLK(clk), .Q(fGy[29]) );
  DFFPOSX1 \fGy_reg[30]  ( .D(n5090), .CLK(clk), .Q(fGy[30]) );
  DFFPOSX1 \Gx_reg[0]  ( .D(n3739), .CLK(clk), .Q(Gx[0]) );
  DFFPOSX1 \Gx_reg[1]  ( .D(n3738), .CLK(clk), .Q(Gx[1]) );
  DFFPOSX1 \fGx_reg[1]  ( .D(n5151), .CLK(clk), .Q(N4390) );
  DFFPOSX1 \Gx_reg[2]  ( .D(n3737), .CLK(clk), .Q(Gx[2]) );
  DFFPOSX1 \fGx_reg[2]  ( .D(n5150), .CLK(clk), .Q(N4387) );
  DFFPOSX1 \Gx_reg[3]  ( .D(n3736), .CLK(clk), .Q(Gx[3]) );
  DFFPOSX1 \fGx_reg[3]  ( .D(n5149), .CLK(clk), .Q(N4384) );
  DFFPOSX1 \Gx_reg[4]  ( .D(n3735), .CLK(clk), .Q(Gx[4]) );
  DFFPOSX1 \fGx_reg[4]  ( .D(n5148), .CLK(clk), .Q(N4381) );
  DFFPOSX1 \Gx_reg[5]  ( .D(n3734), .CLK(clk), .Q(Gx[5]) );
  DFFPOSX1 \fGx_reg[5]  ( .D(n5147), .CLK(clk), .Q(N4378) );
  DFFPOSX1 \Gx_reg[6]  ( .D(n3733), .CLK(clk), .Q(Gx[6]) );
  DFFPOSX1 \fGx_reg[6]  ( .D(n5146), .CLK(clk), .Q(N4375) );
  DFFPOSX1 \Gx_reg[7]  ( .D(n3732), .CLK(clk), .Q(Gx[7]) );
  DFFPOSX1 \fGx_reg[7]  ( .D(n5145), .CLK(clk), .Q(N4372) );
  DFFPOSX1 \Gx_reg[8]  ( .D(n3731), .CLK(clk), .Q(Gx[8]) );
  DFFPOSX1 \fGx_reg[8]  ( .D(n5144), .CLK(clk), .Q(fGx[8]) );
  DFFPOSX1 \Gx_reg[9]  ( .D(n3730), .CLK(clk), .Q(Gx[9]) );
  DFFPOSX1 \fGx_reg[9]  ( .D(n5143), .CLK(clk), .Q(fGx[9]) );
  DFFPOSX1 \Gx_reg[10]  ( .D(n3729), .CLK(clk), .Q(Gx[10]) );
  DFFPOSX1 \fGx_reg[10]  ( .D(n5142), .CLK(clk), .Q(fGx[10]) );
  DFFPOSX1 \Gx_reg[11]  ( .D(n3728), .CLK(clk), .Q(Gx[11]) );
  DFFPOSX1 \fGx_reg[11]  ( .D(n5141), .CLK(clk), .Q(fGx[11]) );
  DFFPOSX1 \Gx_reg[12]  ( .D(n3727), .CLK(clk), .Q(Gx[12]) );
  DFFPOSX1 \fGx_reg[12]  ( .D(n5140), .CLK(clk), .Q(fGx[12]) );
  DFFPOSX1 \Gx_reg[13]  ( .D(n3726), .CLK(clk), .Q(Gx[13]) );
  DFFPOSX1 \fGx_reg[13]  ( .D(n5139), .CLK(clk), .Q(fGx[13]) );
  DFFPOSX1 \Gx_reg[14]  ( .D(n3725), .CLK(clk), .Q(Gx[14]) );
  DFFPOSX1 \fGx_reg[14]  ( .D(n5138), .CLK(clk), .Q(fGx[14]) );
  DFFPOSX1 \Gx_reg[15]  ( .D(n3724), .CLK(clk), .Q(Gx[15]) );
  DFFPOSX1 \fGx_reg[15]  ( .D(n5137), .CLK(clk), .Q(fGx[15]) );
  DFFPOSX1 \Gx_reg[16]  ( .D(n3723), .CLK(clk), .Q(Gx[16]) );
  DFFPOSX1 \fGx_reg[16]  ( .D(n5136), .CLK(clk), .Q(fGx[16]) );
  DFFPOSX1 \Gx_reg[17]  ( .D(n3722), .CLK(clk), .Q(Gx[17]) );
  DFFPOSX1 \fGx_reg[17]  ( .D(n5135), .CLK(clk), .Q(fGx[17]) );
  DFFPOSX1 \Gx_reg[18]  ( .D(n3721), .CLK(clk), .Q(Gx[18]) );
  DFFPOSX1 \fGx_reg[18]  ( .D(n5134), .CLK(clk), .Q(fGx[18]) );
  DFFPOSX1 \Gx_reg[19]  ( .D(n3720), .CLK(clk), .Q(Gx[19]) );
  DFFPOSX1 \fGx_reg[19]  ( .D(n5133), .CLK(clk), .Q(fGx[19]) );
  DFFPOSX1 \Gx_reg[20]  ( .D(n3719), .CLK(clk), .Q(Gx[20]) );
  DFFPOSX1 \fGx_reg[20]  ( .D(n5132), .CLK(clk), .Q(fGx[20]) );
  DFFPOSX1 \Gx_reg[21]  ( .D(n3718), .CLK(clk), .Q(Gx[21]) );
  DFFPOSX1 \fGx_reg[21]  ( .D(n5131), .CLK(clk), .Q(fGx[21]) );
  DFFPOSX1 \Gx_reg[22]  ( .D(n3717), .CLK(clk), .Q(Gx[22]) );
  DFFPOSX1 \fGx_reg[22]  ( .D(n5130), .CLK(clk), .Q(fGx[22]) );
  DFFPOSX1 \Gx_reg[23]  ( .D(n3716), .CLK(clk), .Q(Gx[23]) );
  DFFPOSX1 \fGx_reg[23]  ( .D(n5129), .CLK(clk), .Q(fGx[23]) );
  DFFPOSX1 \Gx_reg[24]  ( .D(n3715), .CLK(clk), .Q(Gx[24]) );
  DFFPOSX1 \fGx_reg[24]  ( .D(n5128), .CLK(clk), .Q(fGx[24]) );
  DFFPOSX1 \Gx_reg[25]  ( .D(n3714), .CLK(clk), .Q(Gx[25]) );
  DFFPOSX1 \fGx_reg[25]  ( .D(n5127), .CLK(clk), .Q(fGx[25]) );
  DFFPOSX1 \Gx_reg[26]  ( .D(n3713), .CLK(clk), .Q(Gx[26]) );
  DFFPOSX1 \fGx_reg[26]  ( .D(n5126), .CLK(clk), .Q(fGx[26]) );
  DFFPOSX1 \Gx_reg[27]  ( .D(n3712), .CLK(clk), .Q(Gx[27]) );
  DFFPOSX1 \fGx_reg[27]  ( .D(n5125), .CLK(clk), .Q(fGx[27]) );
  DFFPOSX1 \Gx_reg[28]  ( .D(n3711), .CLK(clk), .Q(Gx[28]) );
  DFFPOSX1 \fGx_reg[28]  ( .D(n5124), .CLK(clk), .Q(fGx[28]) );
  DFFPOSX1 \Gx_reg[29]  ( .D(n3710), .CLK(clk), .Q(Gx[29]) );
  DFFPOSX1 \fGx_reg[29]  ( .D(n5123), .CLK(clk), .Q(fGx[29]) );
  DFFPOSX1 \Gx_reg[30]  ( .D(n3709), .CLK(clk), .Q(Gx[30]) );
  DFFPOSX1 \fGx_reg[30]  ( .D(n5122), .CLK(clk), .Q(fGx[30]) );
  DFFPOSX1 \Gx_reg[31]  ( .D(n3708), .CLK(clk), .Q(Gx[31]) );
  DFFPOSX1 \fGx_reg[31]  ( .D(n5121), .CLK(clk), .Q(fGx[31]) );
  DFFPOSX1 \fGy_reg[31]  ( .D(n7201), .CLK(clk), .Q(fGy[31]) );
  DFFPOSX1 \tpSum_reg[7]  ( .D(n4660), .CLK(clk), .Q(tpSum[7]) );
  DFFPOSX1 \tpSum_reg[8]  ( .D(n4659), .CLK(clk), .Q(tpSum[8]) );
  DFFPOSX1 \tpSum_reg[9]  ( .D(n4658), .CLK(clk), .Q(tpSum[9]) );
  DFFPOSX1 \tpSum_reg[10]  ( .D(n4657), .CLK(clk), .Q(tpSum[10]) );
  DFFPOSX1 \tpSum_reg[11]  ( .D(n4656), .CLK(clk), .Q(tpSum[11]) );
  DFFPOSX1 \tpSum_reg[12]  ( .D(n4655), .CLK(clk), .Q(tpSum[12]) );
  DFFPOSX1 \tpSum_reg[13]  ( .D(n4654), .CLK(clk), .Q(tpSum[13]) );
  DFFPOSX1 \tpSum_reg[14]  ( .D(n4653), .CLK(clk), .Q(tpSum[14]) );
  DFFPOSX1 \regZ_reg[1][7]  ( .D(n4897), .CLK(clk), .Q(N3796) );
  DFFPOSX1 \regZ_reg[1][6]  ( .D(n4898), .CLK(clk), .Q(N3799) );
  DFFPOSX1 \regZ_reg[1][5]  ( .D(n4899), .CLK(clk), .Q(N3802) );
  DFFPOSX1 \regZ_reg[1][4]  ( .D(n4900), .CLK(clk), .Q(N3805) );
  DFFPOSX1 \regZ_reg[1][3]  ( .D(n4901), .CLK(clk), .Q(N3808) );
  DFFPOSX1 \regZ_reg[1][2]  ( .D(n4902), .CLK(clk), .Q(N3811) );
  DFFPOSX1 \regZ_reg[1][1]  ( .D(n4903), .CLK(clk), .Q(N3814) );
  DFFPOSX1 \regZ_reg[1][0]  ( .D(n4904), .CLK(clk), .Q(N3817) );
  DFFPOSX1 \regZ_tri_enable_reg[1][0]  ( .D(n4704), .CLK(clk), .Q(N3818) );
  DFFPOSX1 \regZ_tri_enable_reg[1][1]  ( .D(n4703), .CLK(clk), .Q(N3815) );
  DFFPOSX1 \regZ_tri_enable_reg[1][2]  ( .D(n4702), .CLK(clk), .Q(N3812) );
  DFFPOSX1 \regZ_tri_enable_reg[1][3]  ( .D(n4701), .CLK(clk), .Q(N3809) );
  DFFPOSX1 \regZ_tri_enable_reg[1][4]  ( .D(n4700), .CLK(clk), .Q(N3806) );
  DFFPOSX1 \regZ_tri_enable_reg[1][5]  ( .D(n4699), .CLK(clk), .Q(N3803) );
  DFFPOSX1 \regZ_tri_enable_reg[1][6]  ( .D(n4698), .CLK(clk), .Q(N3800) );
  DFFPOSX1 \regZ_tri_enable_reg[1][7]  ( .D(n4697), .CLK(clk), .Q(N3797) );
  DFFPOSX1 \regZ_reg[2][7]  ( .D(n4905), .CLK(clk), .Q(N3820) );
  DFFPOSX1 \regZ_reg[2][6]  ( .D(n4906), .CLK(clk), .Q(N3823) );
  DFFPOSX1 \regZ_reg[2][5]  ( .D(n4907), .CLK(clk), .Q(N3826) );
  DFFPOSX1 \regZ_reg[2][4]  ( .D(n4908), .CLK(clk), .Q(N3829) );
  DFFPOSX1 \regZ_reg[2][3]  ( .D(n4909), .CLK(clk), .Q(N3832) );
  DFFPOSX1 \regZ_reg[2][2]  ( .D(n4910), .CLK(clk), .Q(N3835) );
  DFFPOSX1 \regZ_reg[2][1]  ( .D(n4911), .CLK(clk), .Q(N3838) );
  DFFPOSX1 \regZ_reg[2][0]  ( .D(n4912), .CLK(clk), .Q(N3841) );
  DFFPOSX1 \regZ_tri_enable_reg[2][0]  ( .D(n4712), .CLK(clk), .Q(N3842) );
  DFFPOSX1 \regZ_tri_enable_reg[2][1]  ( .D(n4711), .CLK(clk), .Q(N3839) );
  DFFPOSX1 \regZ_tri_enable_reg[2][2]  ( .D(n4710), .CLK(clk), .Q(N3836) );
  DFFPOSX1 \regZ_tri_enable_reg[2][3]  ( .D(n4709), .CLK(clk), .Q(N3833) );
  DFFPOSX1 \regZ_tri_enable_reg[2][4]  ( .D(n4708), .CLK(clk), .Q(N3830) );
  DFFPOSX1 \regZ_tri_enable_reg[2][5]  ( .D(n4707), .CLK(clk), .Q(N3827) );
  DFFPOSX1 \regZ_tri_enable_reg[2][6]  ( .D(n4706), .CLK(clk), .Q(N3824) );
  DFFPOSX1 \regZ_tri_enable_reg[2][7]  ( .D(n4705), .CLK(clk), .Q(N3821) );
  DFFPOSX1 \regZ_reg[10][0]  ( .D(n4976), .CLK(clk), .Q(N4033) );
  DFFPOSX1 \regZ_reg[10][1]  ( .D(n4975), .CLK(clk), .Q(N4030) );
  DFFPOSX1 \regZ_reg[10][2]  ( .D(n4974), .CLK(clk), .Q(N4027) );
  DFFPOSX1 \regZ_reg[10][3]  ( .D(n4973), .CLK(clk), .Q(N4024) );
  DFFPOSX1 \regZ_reg[10][4]  ( .D(n4972), .CLK(clk), .Q(N4021) );
  DFFPOSX1 \regZ_reg[10][5]  ( .D(n4971), .CLK(clk), .Q(N4018) );
  DFFPOSX1 \regZ_reg[10][6]  ( .D(n4970), .CLK(clk), .Q(N4015) );
  DFFPOSX1 \regZ_reg[10][7]  ( .D(n4969), .CLK(clk), .Q(N4012) );
  DFFPOSX1 \regZ_tri_enable_reg[10][7]  ( .D(n4769), .CLK(clk), .Q(N4013) );
  DFFPOSX1 \regZ_tri_enable_reg[10][6]  ( .D(n4770), .CLK(clk), .Q(N4016) );
  DFFPOSX1 \regZ_tri_enable_reg[10][5]  ( .D(n4771), .CLK(clk), .Q(N4019) );
  DFFPOSX1 \regZ_tri_enable_reg[10][4]  ( .D(n4772), .CLK(clk), .Q(N4022) );
  DFFPOSX1 \regZ_tri_enable_reg[10][3]  ( .D(n4773), .CLK(clk), .Q(N4025) );
  DFFPOSX1 \regZ_tri_enable_reg[10][2]  ( .D(n4774), .CLK(clk), .Q(N4028) );
  DFFPOSX1 \regZ_tri_enable_reg[10][1]  ( .D(n4775), .CLK(clk), .Q(N4031) );
  DFFPOSX1 \regZ_tri_enable_reg[10][0]  ( .D(n4776), .CLK(clk), .Q(N4034) );
  DFFPOSX1 \regZ_reg[11][0]  ( .D(n4984), .CLK(clk), .Q(N4057) );
  DFFPOSX1 \regZ_reg[11][1]  ( .D(n4983), .CLK(clk), .Q(N4054) );
  DFFPOSX1 \regZ_reg[11][2]  ( .D(n4982), .CLK(clk), .Q(N4051) );
  DFFPOSX1 \regZ_reg[11][3]  ( .D(n4981), .CLK(clk), .Q(N4048) );
  DFFPOSX1 \regZ_reg[11][4]  ( .D(n4980), .CLK(clk), .Q(N4045) );
  DFFPOSX1 \regZ_reg[11][5]  ( .D(n4979), .CLK(clk), .Q(N4042) );
  DFFPOSX1 \regZ_reg[11][6]  ( .D(n4978), .CLK(clk), .Q(N4039) );
  DFFPOSX1 \regZ_reg[11][7]  ( .D(n4977), .CLK(clk), .Q(N4036) );
  DFFPOSX1 \regZ_tri_enable_reg[11][7]  ( .D(n4777), .CLK(clk), .Q(N4037) );
  DFFPOSX1 \regZ_tri_enable_reg[11][6]  ( .D(n4778), .CLK(clk), .Q(N4040) );
  DFFPOSX1 \regZ_tri_enable_reg[11][5]  ( .D(n4779), .CLK(clk), .Q(N4043) );
  DFFPOSX1 \regZ_tri_enable_reg[11][4]  ( .D(n4780), .CLK(clk), .Q(N4046) );
  DFFPOSX1 \regZ_tri_enable_reg[11][3]  ( .D(n4781), .CLK(clk), .Q(N4049) );
  DFFPOSX1 \regZ_tri_enable_reg[11][2]  ( .D(n4782), .CLK(clk), .Q(N4052) );
  DFFPOSX1 \regZ_tri_enable_reg[11][1]  ( .D(n4783), .CLK(clk), .Q(N4055) );
  DFFPOSX1 \regZ_tri_enable_reg[11][0]  ( .D(n4784), .CLK(clk), .Q(N4058) );
  DFFPOSX1 \regZ_reg[18][0]  ( .D(n5040), .CLK(clk), .Q(N4225) );
  DFFPOSX1 \regZ_reg[18][1]  ( .D(n5039), .CLK(clk), .Q(N4222) );
  DFFPOSX1 \regZ_reg[18][2]  ( .D(n5038), .CLK(clk), .Q(N4219) );
  DFFPOSX1 \regZ_reg[18][3]  ( .D(n5037), .CLK(clk), .Q(N4216) );
  DFFPOSX1 \regZ_reg[18][4]  ( .D(n5036), .CLK(clk), .Q(N4213) );
  DFFPOSX1 \regZ_reg[18][5]  ( .D(n5035), .CLK(clk), .Q(N4210) );
  DFFPOSX1 \regZ_reg[18][6]  ( .D(n5034), .CLK(clk), .Q(N4207) );
  DFFPOSX1 \regZ_reg[18][7]  ( .D(n5033), .CLK(clk), .Q(N4204) );
  DFFPOSX1 \regZ_tri_enable_reg[18][7]  ( .D(n4833), .CLK(clk), .Q(N4205) );
  DFFPOSX1 \regZ_tri_enable_reg[18][6]  ( .D(n4834), .CLK(clk), .Q(N4208) );
  DFFPOSX1 \regZ_tri_enable_reg[18][5]  ( .D(n4835), .CLK(clk), .Q(N4211) );
  DFFPOSX1 \regZ_tri_enable_reg[18][4]  ( .D(n4836), .CLK(clk), .Q(N4214) );
  DFFPOSX1 \regZ_tri_enable_reg[18][3]  ( .D(n4837), .CLK(clk), .Q(N4217) );
  DFFPOSX1 \regZ_tri_enable_reg[18][2]  ( .D(n4838), .CLK(clk), .Q(N4220) );
  DFFPOSX1 \regZ_tri_enable_reg[18][1]  ( .D(n4839), .CLK(clk), .Q(N4223) );
  DFFPOSX1 \regZ_tri_enable_reg[18][0]  ( .D(n4840), .CLK(clk), .Q(N4226) );
  DFFPOSX1 \regZ_reg[19][0]  ( .D(n5048), .CLK(clk), .Q(N4249) );
  DFFPOSX1 \regZ_reg[19][1]  ( .D(n5047), .CLK(clk), .Q(N4246) );
  DFFPOSX1 \regZ_reg[19][2]  ( .D(n5046), .CLK(clk), .Q(N4243) );
  DFFPOSX1 \regZ_reg[19][3]  ( .D(n5045), .CLK(clk), .Q(N4240) );
  DFFPOSX1 \regZ_reg[19][4]  ( .D(n5044), .CLK(clk), .Q(N4237) );
  DFFPOSX1 \regZ_reg[19][5]  ( .D(n5043), .CLK(clk), .Q(N4234) );
  DFFPOSX1 \regZ_reg[19][6]  ( .D(n5042), .CLK(clk), .Q(N4231) );
  DFFPOSX1 \regZ_reg[19][7]  ( .D(n5041), .CLK(clk), .Q(N4228) );
  DFFPOSX1 \regZ_tri_enable_reg[19][7]  ( .D(n4841), .CLK(clk), .Q(N4229) );
  DFFPOSX1 \regZ_tri_enable_reg[19][6]  ( .D(n4842), .CLK(clk), .Q(N4232) );
  DFFPOSX1 \regZ_tri_enable_reg[19][5]  ( .D(n4843), .CLK(clk), .Q(N4235) );
  DFFPOSX1 \regZ_tri_enable_reg[19][4]  ( .D(n4844), .CLK(clk), .Q(N4238) );
  DFFPOSX1 \regZ_tri_enable_reg[19][3]  ( .D(n4845), .CLK(clk), .Q(N4241) );
  DFFPOSX1 \regZ_tri_enable_reg[19][2]  ( .D(n4846), .CLK(clk), .Q(N4244) );
  DFFPOSX1 \regZ_tri_enable_reg[19][1]  ( .D(n4847), .CLK(clk), .Q(N4247) );
  DFFPOSX1 \regZ_tri_enable_reg[19][0]  ( .D(n4848), .CLK(clk), .Q(N4250) );
  DFFPOSX1 \regZ_reg[12][0]  ( .D(n4985), .CLK(clk), .Q(N4081) );
  DFFPOSX1 \regZ_reg[12][7]  ( .D(n4986), .CLK(clk), .Q(N4060) );
  DFFPOSX1 \regZ_reg[12][6]  ( .D(n4987), .CLK(clk), .Q(N4063) );
  DFFPOSX1 \regZ_reg[12][5]  ( .D(n4988), .CLK(clk), .Q(N4066) );
  DFFPOSX1 \regZ_reg[12][4]  ( .D(n4989), .CLK(clk), .Q(N4069) );
  DFFPOSX1 \regZ_reg[12][3]  ( .D(n4990), .CLK(clk), .Q(N4072) );
  DFFPOSX1 \regZ_reg[12][2]  ( .D(n4991), .CLK(clk), .Q(N4075) );
  DFFPOSX1 \regZ_reg[12][1]  ( .D(n4992), .CLK(clk), .Q(N4078) );
  DFFPOSX1 \regZ_tri_enable_reg[12][0]  ( .D(n4792), .CLK(clk), .Q(N4082) );
  DFFPOSX1 \regZ_tri_enable_reg[12][1]  ( .D(n4791), .CLK(clk), .Q(N4079) );
  DFFPOSX1 \regZ_tri_enable_reg[12][2]  ( .D(n4790), .CLK(clk), .Q(N4076) );
  DFFPOSX1 \regZ_tri_enable_reg[12][3]  ( .D(n4789), .CLK(clk), .Q(N4073) );
  DFFPOSX1 \regZ_tri_enable_reg[12][4]  ( .D(n4788), .CLK(clk), .Q(N4070) );
  DFFPOSX1 \regZ_tri_enable_reg[12][5]  ( .D(n4787), .CLK(clk), .Q(N4067) );
  DFFPOSX1 \regZ_tri_enable_reg[12][6]  ( .D(n4786), .CLK(clk), .Q(N4064) );
  DFFPOSX1 \regZ_tri_enable_reg[12][7]  ( .D(n4785), .CLK(clk), .Q(N4061) );
  DFFPOSX1 \regZ_reg[13][0]  ( .D(n5000), .CLK(clk), .Q(N4105) );
  DFFPOSX1 \regZ_reg[13][1]  ( .D(n4999), .CLK(clk), .Q(N4102) );
  DFFPOSX1 \regZ_reg[13][2]  ( .D(n4998), .CLK(clk), .Q(N4099) );
  DFFPOSX1 \regZ_reg[13][3]  ( .D(n4997), .CLK(clk), .Q(N4096) );
  DFFPOSX1 \regZ_reg[13][4]  ( .D(n4996), .CLK(clk), .Q(N4093) );
  DFFPOSX1 \regZ_reg[13][5]  ( .D(n4995), .CLK(clk), .Q(N4090) );
  DFFPOSX1 \regZ_reg[13][6]  ( .D(n4994), .CLK(clk), .Q(N4087) );
  DFFPOSX1 \regZ_reg[13][7]  ( .D(n4993), .CLK(clk), .Q(N4084) );
  DFFPOSX1 \regZ_tri_enable_reg[13][7]  ( .D(n4793), .CLK(clk), .Q(N4085) );
  DFFPOSX1 \regZ_tri_enable_reg[13][6]  ( .D(n4794), .CLK(clk), .Q(N4088) );
  DFFPOSX1 \regZ_tri_enable_reg[13][5]  ( .D(n4795), .CLK(clk), .Q(N4091) );
  DFFPOSX1 \regZ_tri_enable_reg[13][4]  ( .D(n4796), .CLK(clk), .Q(N4094) );
  DFFPOSX1 \regZ_tri_enable_reg[13][3]  ( .D(n4797), .CLK(clk), .Q(N4097) );
  DFFPOSX1 \regZ_tri_enable_reg[13][2]  ( .D(n4798), .CLK(clk), .Q(N4100) );
  DFFPOSX1 \regZ_tri_enable_reg[13][1]  ( .D(n4799), .CLK(clk), .Q(N4103) );
  DFFPOSX1 \regZ_tri_enable_reg[13][0]  ( .D(n4800), .CLK(clk), .Q(N4106) );
  DFFPOSX1 \regZ_reg[20][0]  ( .D(n5056), .CLK(clk), .Q(N4273) );
  DFFPOSX1 \regZ_reg[20][1]  ( .D(n5055), .CLK(clk), .Q(N4270) );
  DFFPOSX1 \regZ_reg[20][2]  ( .D(n5054), .CLK(clk), .Q(N4267) );
  DFFPOSX1 \regZ_reg[20][3]  ( .D(n5053), .CLK(clk), .Q(N4264) );
  DFFPOSX1 \regZ_reg[20][4]  ( .D(n5052), .CLK(clk), .Q(N4261) );
  DFFPOSX1 \regZ_reg[20][5]  ( .D(n5051), .CLK(clk), .Q(N4258) );
  DFFPOSX1 \regZ_reg[20][6]  ( .D(n5050), .CLK(clk), .Q(N4255) );
  DFFPOSX1 \regZ_reg[20][7]  ( .D(n5049), .CLK(clk), .Q(N4252) );
  DFFPOSX1 \regZ_tri_enable_reg[20][7]  ( .D(n4849), .CLK(clk), .Q(N4253) );
  DFFPOSX1 \regZ_tri_enable_reg[20][6]  ( .D(n4850), .CLK(clk), .Q(N4256) );
  DFFPOSX1 \regZ_tri_enable_reg[20][5]  ( .D(n4851), .CLK(clk), .Q(N4259) );
  DFFPOSX1 \regZ_tri_enable_reg[20][4]  ( .D(n4852), .CLK(clk), .Q(N4262) );
  DFFPOSX1 \regZ_tri_enable_reg[20][3]  ( .D(n4853), .CLK(clk), .Q(N4265) );
  DFFPOSX1 \regZ_tri_enable_reg[20][2]  ( .D(n4854), .CLK(clk), .Q(N4268) );
  DFFPOSX1 \regZ_tri_enable_reg[20][1]  ( .D(n4855), .CLK(clk), .Q(N4271) );
  DFFPOSX1 \regZ_tri_enable_reg[20][0]  ( .D(n4856), .CLK(clk), .Q(N4274) );
  DFFPOSX1 \regZ_reg[21][0]  ( .D(n5064), .CLK(clk), .Q(N4297) );
  DFFPOSX1 \regZ_reg[21][1]  ( .D(n5063), .CLK(clk), .Q(N4294) );
  DFFPOSX1 \regZ_reg[21][2]  ( .D(n5062), .CLK(clk), .Q(N4291) );
  DFFPOSX1 \regZ_reg[21][3]  ( .D(n5061), .CLK(clk), .Q(N4288) );
  DFFPOSX1 \regZ_reg[21][4]  ( .D(n5060), .CLK(clk), .Q(N4285) );
  DFFPOSX1 \regZ_reg[21][5]  ( .D(n5059), .CLK(clk), .Q(N4282) );
  DFFPOSX1 \regZ_reg[21][6]  ( .D(n5058), .CLK(clk), .Q(N4279) );
  DFFPOSX1 \regZ_reg[21][7]  ( .D(n5057), .CLK(clk), .Q(N4276) );
  DFFPOSX1 \regZ_tri_enable_reg[21][7]  ( .D(n4857), .CLK(clk), .Q(N4277) );
  DFFPOSX1 \regZ_tri_enable_reg[21][6]  ( .D(n4858), .CLK(clk), .Q(N4280) );
  DFFPOSX1 \regZ_tri_enable_reg[21][5]  ( .D(n4859), .CLK(clk), .Q(N4283) );
  DFFPOSX1 \regZ_tri_enable_reg[21][4]  ( .D(n4860), .CLK(clk), .Q(N4286) );
  DFFPOSX1 \regZ_tri_enable_reg[21][3]  ( .D(n4861), .CLK(clk), .Q(N4289) );
  DFFPOSX1 \regZ_tri_enable_reg[21][2]  ( .D(n4862), .CLK(clk), .Q(N4292) );
  DFFPOSX1 \regZ_tri_enable_reg[21][1]  ( .D(n4863), .CLK(clk), .Q(N4295) );
  DFFPOSX1 \regZ_tri_enable_reg[21][0]  ( .D(n4864), .CLK(clk), .Q(N4298) );
  DFFPOSX1 \regZ_reg[14][0]  ( .D(n5008), .CLK(clk), .Q(N4129) );
  DFFPOSX1 \regZ_reg[14][1]  ( .D(n5007), .CLK(clk), .Q(N4126) );
  DFFPOSX1 \regZ_reg[14][2]  ( .D(n5006), .CLK(clk), .Q(N4123) );
  DFFPOSX1 \regZ_reg[14][3]  ( .D(n5005), .CLK(clk), .Q(N4120) );
  DFFPOSX1 \regZ_reg[14][4]  ( .D(n5004), .CLK(clk), .Q(N4117) );
  DFFPOSX1 \regZ_reg[14][5]  ( .D(n5003), .CLK(clk), .Q(N4114) );
  DFFPOSX1 \regZ_reg[14][6]  ( .D(n5002), .CLK(clk), .Q(N4111) );
  DFFPOSX1 \regZ_reg[14][7]  ( .D(n5001), .CLK(clk), .Q(N4108) );
  DFFPOSX1 \regZ_tri_enable_reg[14][7]  ( .D(n4801), .CLK(clk), .Q(N4109) );
  DFFPOSX1 \regZ_tri_enable_reg[14][6]  ( .D(n4802), .CLK(clk), .Q(N4112) );
  DFFPOSX1 \regZ_tri_enable_reg[14][5]  ( .D(n4803), .CLK(clk), .Q(N4115) );
  DFFPOSX1 \regZ_tri_enable_reg[14][4]  ( .D(n4804), .CLK(clk), .Q(N4118) );
  DFFPOSX1 \regZ_tri_enable_reg[14][3]  ( .D(n4805), .CLK(clk), .Q(N4121) );
  DFFPOSX1 \regZ_tri_enable_reg[14][2]  ( .D(n4806), .CLK(clk), .Q(N4124) );
  DFFPOSX1 \regZ_tri_enable_reg[14][1]  ( .D(n4807), .CLK(clk), .Q(N4127) );
  DFFPOSX1 \regZ_tri_enable_reg[14][0]  ( .D(n4808), .CLK(clk), .Q(N4130) );
  DFFPOSX1 \regZ_reg[15][0]  ( .D(n5016), .CLK(clk), .Q(N4153) );
  DFFPOSX1 \regZ_reg[15][1]  ( .D(n5015), .CLK(clk), .Q(N4150) );
  DFFPOSX1 \regZ_reg[15][2]  ( .D(n5014), .CLK(clk), .Q(N4147) );
  DFFPOSX1 \regZ_reg[15][3]  ( .D(n5013), .CLK(clk), .Q(N4144) );
  DFFPOSX1 \regZ_reg[15][4]  ( .D(n5012), .CLK(clk), .Q(N4141) );
  DFFPOSX1 \regZ_reg[15][5]  ( .D(n5011), .CLK(clk), .Q(N4138) );
  DFFPOSX1 \regZ_reg[15][6]  ( .D(n5010), .CLK(clk), .Q(N4135) );
  DFFPOSX1 \regZ_reg[15][7]  ( .D(n5009), .CLK(clk), .Q(N4132) );
  DFFPOSX1 \regZ_tri_enable_reg[15][7]  ( .D(n4809), .CLK(clk), .Q(N4133) );
  DFFPOSX1 \regZ_tri_enable_reg[15][6]  ( .D(n4810), .CLK(clk), .Q(N4136) );
  DFFPOSX1 \regZ_tri_enable_reg[15][5]  ( .D(n4811), .CLK(clk), .Q(N4139) );
  DFFPOSX1 \regZ_tri_enable_reg[15][4]  ( .D(n4812), .CLK(clk), .Q(N4142) );
  DFFPOSX1 \regZ_tri_enable_reg[15][3]  ( .D(n4813), .CLK(clk), .Q(N4145) );
  DFFPOSX1 \regZ_tri_enable_reg[15][2]  ( .D(n4814), .CLK(clk), .Q(N4148) );
  DFFPOSX1 \regZ_tri_enable_reg[15][1]  ( .D(n4815), .CLK(clk), .Q(N4151) );
  DFFPOSX1 \regZ_tri_enable_reg[15][0]  ( .D(n4816), .CLK(clk), .Q(N4154) );
  DFFPOSX1 \regZ_reg[22][0]  ( .D(n5072), .CLK(clk), .Q(N4321) );
  DFFPOSX1 \regZ_reg[22][1]  ( .D(n5071), .CLK(clk), .Q(N4318) );
  DFFPOSX1 \regZ_reg[22][2]  ( .D(n5070), .CLK(clk), .Q(N4315) );
  DFFPOSX1 \regZ_reg[22][3]  ( .D(n5069), .CLK(clk), .Q(N4312) );
  DFFPOSX1 \regZ_reg[22][4]  ( .D(n5068), .CLK(clk), .Q(N4309) );
  DFFPOSX1 \regZ_reg[22][5]  ( .D(n5067), .CLK(clk), .Q(N4306) );
  DFFPOSX1 \regZ_reg[22][6]  ( .D(n5066), .CLK(clk), .Q(N4303) );
  DFFPOSX1 \regZ_reg[22][7]  ( .D(n5065), .CLK(clk), .Q(N4300) );
  DFFPOSX1 \regZ_tri_enable_reg[22][7]  ( .D(n4865), .CLK(clk), .Q(N4301) );
  DFFPOSX1 \regZ_tri_enable_reg[22][6]  ( .D(n4866), .CLK(clk), .Q(N4304) );
  DFFPOSX1 \regZ_tri_enable_reg[22][5]  ( .D(n4867), .CLK(clk), .Q(N4307) );
  DFFPOSX1 \regZ_tri_enable_reg[22][4]  ( .D(n4868), .CLK(clk), .Q(N4310) );
  DFFPOSX1 \regZ_tri_enable_reg[22][3]  ( .D(n4869), .CLK(clk), .Q(N4313) );
  DFFPOSX1 \regZ_tri_enable_reg[22][2]  ( .D(n4870), .CLK(clk), .Q(N4316) );
  DFFPOSX1 \regZ_tri_enable_reg[22][1]  ( .D(n4871), .CLK(clk), .Q(N4319) );
  DFFPOSX1 \regZ_tri_enable_reg[22][0]  ( .D(n4872), .CLK(clk), .Q(N4322) );
  DFFPOSX1 \regZ_reg[23][0]  ( .D(n5080), .CLK(clk), .Q(N4345) );
  DFFPOSX1 \regZ_reg[23][1]  ( .D(n5079), .CLK(clk), .Q(N4342) );
  DFFPOSX1 \regZ_reg[23][2]  ( .D(n5078), .CLK(clk), .Q(N4339) );
  DFFPOSX1 \regZ_reg[23][3]  ( .D(n5077), .CLK(clk), .Q(N4336) );
  DFFPOSX1 \regZ_reg[23][4]  ( .D(n5076), .CLK(clk), .Q(N4333) );
  DFFPOSX1 \regZ_reg[23][5]  ( .D(n5075), .CLK(clk), .Q(N4330) );
  DFFPOSX1 \regZ_reg[23][6]  ( .D(n5074), .CLK(clk), .Q(N4327) );
  DFFPOSX1 \regZ_reg[23][7]  ( .D(n5073), .CLK(clk), .Q(N4324) );
  DFFPOSX1 \regZ_tri_enable_reg[23][7]  ( .D(n4873), .CLK(clk), .Q(N4325) );
  DFFPOSX1 \regZ_tri_enable_reg[23][6]  ( .D(n4874), .CLK(clk), .Q(N4328) );
  DFFPOSX1 \regZ_tri_enable_reg[23][5]  ( .D(n4875), .CLK(clk), .Q(N4331) );
  DFFPOSX1 \regZ_tri_enable_reg[23][4]  ( .D(n4876), .CLK(clk), .Q(N4334) );
  DFFPOSX1 \regZ_tri_enable_reg[23][3]  ( .D(n4877), .CLK(clk), .Q(N4337) );
  DFFPOSX1 \regZ_tri_enable_reg[23][2]  ( .D(n4878), .CLK(clk), .Q(N4340) );
  DFFPOSX1 \regZ_tri_enable_reg[23][1]  ( .D(n4879), .CLK(clk), .Q(N4343) );
  DFFPOSX1 \regZ_tri_enable_reg[23][0]  ( .D(n4880), .CLK(clk), .Q(N4346) );
  DFFPOSX1 \regZ_reg[24][7]  ( .D(n5081), .CLK(clk), .Q(N4348) );
  DFFPOSX1 \regZ_reg[24][6]  ( .D(n5082), .CLK(clk), .Q(N4351) );
  DFFPOSX1 \regZ_reg[24][5]  ( .D(n5083), .CLK(clk), .Q(N4354) );
  DFFPOSX1 \regZ_reg[24][4]  ( .D(n5084), .CLK(clk), .Q(N4357) );
  DFFPOSX1 \regZ_reg[24][3]  ( .D(n5085), .CLK(clk), .Q(N4360) );
  DFFPOSX1 \regZ_reg[24][2]  ( .D(n5086), .CLK(clk), .Q(N4363) );
  DFFPOSX1 \regZ_reg[24][1]  ( .D(n5087), .CLK(clk), .Q(N4366) );
  DFFPOSX1 \regZ_reg[24][0]  ( .D(n5088), .CLK(clk), .Q(N4369) );
  DFFPOSX1 \regZ_tri_enable_reg[24][0]  ( .D(n4888), .CLK(clk), .Q(N4370) );
  DFFPOSX1 \regZ_tri_enable_reg[24][1]  ( .D(n4887), .CLK(clk), .Q(N4367) );
  DFFPOSX1 \regZ_tri_enable_reg[24][2]  ( .D(n4886), .CLK(clk), .Q(N4364) );
  DFFPOSX1 \regZ_tri_enable_reg[24][3]  ( .D(n4885), .CLK(clk), .Q(N4361) );
  DFFPOSX1 \regZ_tri_enable_reg[24][4]  ( .D(n4884), .CLK(clk), .Q(N4358) );
  DFFPOSX1 \regZ_tri_enable_reg[24][5]  ( .D(n4883), .CLK(clk), .Q(N4355) );
  DFFPOSX1 \regZ_tri_enable_reg[24][6]  ( .D(n4882), .CLK(clk), .Q(N4352) );
  DFFPOSX1 \regZ_tri_enable_reg[24][7]  ( .D(n4881), .CLK(clk), .Q(N4349) );
  DFFPOSX1 \regZ_reg[17][7]  ( .D(n5025), .CLK(clk), .Q(N4180) );
  DFFPOSX1 \regZ_reg[17][6]  ( .D(n5026), .CLK(clk), .Q(N4183) );
  DFFPOSX1 \regZ_reg[17][5]  ( .D(n5027), .CLK(clk), .Q(N4186) );
  DFFPOSX1 \regZ_reg[17][4]  ( .D(n5028), .CLK(clk), .Q(N4189) );
  DFFPOSX1 \regZ_reg[17][3]  ( .D(n5029), .CLK(clk), .Q(N4192) );
  DFFPOSX1 \regZ_reg[17][2]  ( .D(n5030), .CLK(clk), .Q(N4195) );
  DFFPOSX1 \regZ_reg[17][1]  ( .D(n5031), .CLK(clk), .Q(N4198) );
  DFFPOSX1 \regZ_reg[17][0]  ( .D(n5032), .CLK(clk), .Q(N4201) );
  DFFPOSX1 \regZ_tri_enable_reg[17][0]  ( .D(n4832), .CLK(clk), .Q(N4202) );
  DFFPOSX1 \regZ_tri_enable_reg[17][1]  ( .D(n4831), .CLK(clk), .Q(N4199) );
  DFFPOSX1 \regZ_tri_enable_reg[17][2]  ( .D(n4830), .CLK(clk), .Q(N4196) );
  DFFPOSX1 \regZ_tri_enable_reg[17][3]  ( .D(n4829), .CLK(clk), .Q(N4193) );
  DFFPOSX1 \regZ_tri_enable_reg[17][4]  ( .D(n4828), .CLK(clk), .Q(N4190) );
  DFFPOSX1 \regZ_tri_enable_reg[17][5]  ( .D(n4827), .CLK(clk), .Q(N4187) );
  DFFPOSX1 \regZ_tri_enable_reg[17][6]  ( .D(n4826), .CLK(clk), .Q(N4184) );
  DFFPOSX1 \regZ_tri_enable_reg[17][7]  ( .D(n4825), .CLK(clk), .Q(N4181) );
  DFFPOSX1 \regZ_reg[16][7]  ( .D(n5017), .CLK(clk), .Q(N4156) );
  DFFPOSX1 \regZ_reg[16][6]  ( .D(n5018), .CLK(clk), .Q(N4159) );
  DFFPOSX1 \regZ_reg[16][5]  ( .D(n5019), .CLK(clk), .Q(N4162) );
  DFFPOSX1 \regZ_reg[16][4]  ( .D(n5020), .CLK(clk), .Q(N4165) );
  DFFPOSX1 \regZ_reg[16][3]  ( .D(n5021), .CLK(clk), .Q(N4168) );
  DFFPOSX1 \regZ_reg[16][2]  ( .D(n5022), .CLK(clk), .Q(N4171) );
  DFFPOSX1 \regZ_reg[16][1]  ( .D(n5023), .CLK(clk), .Q(N4174) );
  DFFPOSX1 \regZ_reg[16][0]  ( .D(n5024), .CLK(clk), .Q(N4177) );
  DFFPOSX1 \regZ_tri_enable_reg[16][0]  ( .D(n4824), .CLK(clk), .Q(N4178) );
  DFFPOSX1 \regZ_tri_enable_reg[16][1]  ( .D(n4823), .CLK(clk), .Q(N4175) );
  DFFPOSX1 \regZ_tri_enable_reg[16][2]  ( .D(n4822), .CLK(clk), .Q(N4172) );
  DFFPOSX1 \regZ_tri_enable_reg[16][3]  ( .D(n4821), .CLK(clk), .Q(N4169) );
  DFFPOSX1 \regZ_tri_enable_reg[16][4]  ( .D(n4820), .CLK(clk), .Q(N4166) );
  DFFPOSX1 \regZ_tri_enable_reg[16][5]  ( .D(n4819), .CLK(clk), .Q(N4163) );
  DFFPOSX1 \regZ_tri_enable_reg[16][6]  ( .D(n4818), .CLK(clk), .Q(N4160) );
  DFFPOSX1 \regZ_tri_enable_reg[16][7]  ( .D(n4817), .CLK(clk), .Q(N4157) );
  DFFPOSX1 \regZ_reg[9][7]  ( .D(n4961), .CLK(clk), .Q(N3988) );
  DFFPOSX1 \regZ_reg[9][6]  ( .D(n4962), .CLK(clk), .Q(N3991) );
  DFFPOSX1 \regZ_reg[9][5]  ( .D(n4963), .CLK(clk), .Q(N3994) );
  DFFPOSX1 \regZ_reg[9][4]  ( .D(n4964), .CLK(clk), .Q(N3997) );
  DFFPOSX1 \regZ_reg[9][3]  ( .D(n4965), .CLK(clk), .Q(N4000) );
  DFFPOSX1 \regZ_reg[9][2]  ( .D(n4966), .CLK(clk), .Q(N4003) );
  DFFPOSX1 \regZ_reg[9][1]  ( .D(n4967), .CLK(clk), .Q(N4006) );
  DFFPOSX1 \regZ_reg[9][0]  ( .D(n4968), .CLK(clk), .Q(N4009) );
  DFFPOSX1 \regZ_tri_enable_reg[9][0]  ( .D(n4768), .CLK(clk), .Q(N4010) );
  DFFPOSX1 \regZ_tri_enable_reg[9][1]  ( .D(n4767), .CLK(clk), .Q(N4007) );
  DFFPOSX1 \regZ_tri_enable_reg[9][2]  ( .D(n4766), .CLK(clk), .Q(N4004) );
  DFFPOSX1 \regZ_tri_enable_reg[9][3]  ( .D(n4765), .CLK(clk), .Q(N4001) );
  DFFPOSX1 \regZ_tri_enable_reg[9][4]  ( .D(n4764), .CLK(clk), .Q(N3998) );
  DFFPOSX1 \regZ_tri_enable_reg[9][5]  ( .D(n4763), .CLK(clk), .Q(N3995) );
  DFFPOSX1 \regZ_tri_enable_reg[9][6]  ( .D(n4762), .CLK(clk), .Q(N3992) );
  DFFPOSX1 \regZ_tri_enable_reg[9][7]  ( .D(n4761), .CLK(clk), .Q(N3989) );
  DFFPOSX1 \regZ_reg[8][7]  ( .D(n4953), .CLK(clk), .Q(N3964) );
  DFFPOSX1 \regZ_reg[8][6]  ( .D(n4954), .CLK(clk), .Q(N3967) );
  DFFPOSX1 \regZ_reg[8][5]  ( .D(n4955), .CLK(clk), .Q(N3970) );
  DFFPOSX1 \regZ_reg[8][4]  ( .D(n4956), .CLK(clk), .Q(N3973) );
  DFFPOSX1 \regZ_reg[8][3]  ( .D(n4957), .CLK(clk), .Q(N3976) );
  DFFPOSX1 \regZ_reg[8][2]  ( .D(n4958), .CLK(clk), .Q(N3979) );
  DFFPOSX1 \regZ_reg[8][1]  ( .D(n4959), .CLK(clk), .Q(N3982) );
  DFFPOSX1 \regZ_reg[8][0]  ( .D(n4960), .CLK(clk), .Q(N3985) );
  DFFPOSX1 \regZ_tri_enable_reg[8][0]  ( .D(n4760), .CLK(clk), .Q(N3986) );
  DFFPOSX1 \regZ_tri_enable_reg[8][1]  ( .D(n4759), .CLK(clk), .Q(N3983) );
  DFFPOSX1 \regZ_tri_enable_reg[8][2]  ( .D(n4758), .CLK(clk), .Q(N3980) );
  DFFPOSX1 \regZ_tri_enable_reg[8][3]  ( .D(n4757), .CLK(clk), .Q(N3977) );
  DFFPOSX1 \regZ_tri_enable_reg[8][4]  ( .D(n4756), .CLK(clk), .Q(N3974) );
  DFFPOSX1 \regZ_tri_enable_reg[8][5]  ( .D(n4755), .CLK(clk), .Q(N3971) );
  DFFPOSX1 \regZ_tri_enable_reg[8][6]  ( .D(n4754), .CLK(clk), .Q(N3968) );
  DFFPOSX1 \regZ_tri_enable_reg[8][7]  ( .D(n4753), .CLK(clk), .Q(N3965) );
  DFFPOSX1 \regZ_reg[7][7]  ( .D(n4945), .CLK(clk), .Q(N3940) );
  DFFPOSX1 \regZ_reg[7][6]  ( .D(n4946), .CLK(clk), .Q(N3943) );
  DFFPOSX1 \regZ_reg[7][5]  ( .D(n4947), .CLK(clk), .Q(N3946) );
  DFFPOSX1 \regZ_reg[7][4]  ( .D(n4948), .CLK(clk), .Q(N3949) );
  DFFPOSX1 \regZ_reg[7][3]  ( .D(n4949), .CLK(clk), .Q(N3952) );
  DFFPOSX1 \regZ_reg[7][2]  ( .D(n4950), .CLK(clk), .Q(N3955) );
  DFFPOSX1 \regZ_reg[7][1]  ( .D(n4951), .CLK(clk), .Q(N3958) );
  DFFPOSX1 \regZ_reg[7][0]  ( .D(n4952), .CLK(clk), .Q(N3961) );
  DFFPOSX1 \regZ_tri_enable_reg[7][0]  ( .D(n4752), .CLK(clk), .Q(N3962) );
  DFFPOSX1 \regZ_tri_enable_reg[7][1]  ( .D(n4751), .CLK(clk), .Q(N3959) );
  DFFPOSX1 \regZ_tri_enable_reg[7][2]  ( .D(n4750), .CLK(clk), .Q(N3956) );
  DFFPOSX1 \regZ_tri_enable_reg[7][3]  ( .D(n4749), .CLK(clk), .Q(N3953) );
  DFFPOSX1 \regZ_tri_enable_reg[7][4]  ( .D(n4748), .CLK(clk), .Q(N3950) );
  DFFPOSX1 \regZ_tri_enable_reg[7][5]  ( .D(n4747), .CLK(clk), .Q(N3947) );
  DFFPOSX1 \regZ_tri_enable_reg[7][6]  ( .D(n4746), .CLK(clk), .Q(N3944) );
  DFFPOSX1 \regZ_tri_enable_reg[7][7]  ( .D(n4745), .CLK(clk), .Q(N3941) );
  DFFPOSX1 \regZ_reg[6][7]  ( .D(n4937), .CLK(clk), .Q(N3916) );
  DFFPOSX1 \regZ_reg[6][6]  ( .D(n4938), .CLK(clk), .Q(N3919) );
  DFFPOSX1 \regZ_reg[6][5]  ( .D(n4939), .CLK(clk), .Q(N3922) );
  DFFPOSX1 \regZ_reg[6][4]  ( .D(n4940), .CLK(clk), .Q(N3925) );
  DFFPOSX1 \regZ_reg[6][3]  ( .D(n4941), .CLK(clk), .Q(N3928) );
  DFFPOSX1 \regZ_reg[6][2]  ( .D(n4942), .CLK(clk), .Q(N3931) );
  DFFPOSX1 \regZ_reg[6][1]  ( .D(n4943), .CLK(clk), .Q(N3934) );
  DFFPOSX1 \regZ_reg[6][0]  ( .D(n4944), .CLK(clk), .Q(N3937) );
  DFFPOSX1 \regZ_tri_enable_reg[6][0]  ( .D(n4744), .CLK(clk), .Q(N3938) );
  DFFPOSX1 \regZ_tri_enable_reg[6][1]  ( .D(n4743), .CLK(clk), .Q(N3935) );
  DFFPOSX1 \regZ_tri_enable_reg[6][2]  ( .D(n4742), .CLK(clk), .Q(N3932) );
  DFFPOSX1 \regZ_tri_enable_reg[6][3]  ( .D(n4741), .CLK(clk), .Q(N3929) );
  DFFPOSX1 \regZ_tri_enable_reg[6][4]  ( .D(n4740), .CLK(clk), .Q(N3926) );
  DFFPOSX1 \regZ_tri_enable_reg[6][5]  ( .D(n4739), .CLK(clk), .Q(N3923) );
  DFFPOSX1 \regZ_tri_enable_reg[6][6]  ( .D(n4738), .CLK(clk), .Q(N3920) );
  DFFPOSX1 \regZ_tri_enable_reg[6][7]  ( .D(n4737), .CLK(clk), .Q(N3917) );
  DFFPOSX1 \regZ_reg[5][7]  ( .D(n4929), .CLK(clk), .Q(N3892) );
  DFFPOSX1 \regZ_reg[5][6]  ( .D(n4930), .CLK(clk), .Q(N3895) );
  DFFPOSX1 \regZ_reg[5][5]  ( .D(n4931), .CLK(clk), .Q(N3898) );
  DFFPOSX1 \regZ_reg[5][4]  ( .D(n4932), .CLK(clk), .Q(N3901) );
  DFFPOSX1 \regZ_reg[5][3]  ( .D(n4933), .CLK(clk), .Q(N3904) );
  DFFPOSX1 \regZ_reg[5][2]  ( .D(n4934), .CLK(clk), .Q(N3907) );
  DFFPOSX1 \regZ_reg[5][1]  ( .D(n4935), .CLK(clk), .Q(N3910) );
  DFFPOSX1 \regZ_reg[5][0]  ( .D(n4936), .CLK(clk), .Q(N3913) );
  DFFPOSX1 \regZ_tri_enable_reg[5][0]  ( .D(n4736), .CLK(clk), .Q(N3914) );
  DFFPOSX1 \regZ_tri_enable_reg[5][1]  ( .D(n4735), .CLK(clk), .Q(N3911) );
  DFFPOSX1 \regZ_tri_enable_reg[5][2]  ( .D(n4734), .CLK(clk), .Q(N3908) );
  DFFPOSX1 \regZ_tri_enable_reg[5][3]  ( .D(n4733), .CLK(clk), .Q(N3905) );
  DFFPOSX1 \regZ_tri_enable_reg[5][4]  ( .D(n4732), .CLK(clk), .Q(N3902) );
  DFFPOSX1 \regZ_tri_enable_reg[5][5]  ( .D(n4731), .CLK(clk), .Q(N3899) );
  DFFPOSX1 \regZ_tri_enable_reg[5][6]  ( .D(n4730), .CLK(clk), .Q(N3896) );
  DFFPOSX1 \regZ_tri_enable_reg[5][7]  ( .D(n4729), .CLK(clk), .Q(N3893) );
  DFFPOSX1 \regZ_reg[4][7]  ( .D(n4921), .CLK(clk), .Q(N3868) );
  DFFPOSX1 \regZ_reg[4][6]  ( .D(n4922), .CLK(clk), .Q(N3871) );
  DFFPOSX1 \regZ_reg[4][5]  ( .D(n4923), .CLK(clk), .Q(N3874) );
  DFFPOSX1 \regZ_reg[4][4]  ( .D(n4924), .CLK(clk), .Q(N3877) );
  DFFPOSX1 \regZ_reg[4][3]  ( .D(n4925), .CLK(clk), .Q(N3880) );
  DFFPOSX1 \regZ_reg[4][2]  ( .D(n4926), .CLK(clk), .Q(N3883) );
  DFFPOSX1 \regZ_reg[4][1]  ( .D(n4927), .CLK(clk), .Q(N3886) );
  DFFPOSX1 \regZ_reg[4][0]  ( .D(n4928), .CLK(clk), .Q(N3889) );
  DFFPOSX1 \regZ_tri_enable_reg[4][0]  ( .D(n4728), .CLK(clk), .Q(N3890) );
  DFFPOSX1 \regZ_tri_enable_reg[4][1]  ( .D(n4727), .CLK(clk), .Q(N3887) );
  DFFPOSX1 \regZ_tri_enable_reg[4][2]  ( .D(n4726), .CLK(clk), .Q(N3884) );
  DFFPOSX1 \regZ_tri_enable_reg[4][3]  ( .D(n4725), .CLK(clk), .Q(N3881) );
  DFFPOSX1 \regZ_tri_enable_reg[4][4]  ( .D(n4724), .CLK(clk), .Q(N3878) );
  DFFPOSX1 \regZ_tri_enable_reg[4][5]  ( .D(n4723), .CLK(clk), .Q(N3875) );
  DFFPOSX1 \regZ_tri_enable_reg[4][6]  ( .D(n4722), .CLK(clk), .Q(N3872) );
  DFFPOSX1 \regZ_tri_enable_reg[4][7]  ( .D(n4721), .CLK(clk), .Q(N3869) );
  DFFPOSX1 \regZ_reg[3][7]  ( .D(n4913), .CLK(clk), .Q(N3844) );
  DFFPOSX1 \regZ_reg[3][6]  ( .D(n4914), .CLK(clk), .Q(N3847) );
  DFFPOSX1 \regZ_reg[3][5]  ( .D(n4915), .CLK(clk), .Q(N3850) );
  DFFPOSX1 \regZ_reg[3][4]  ( .D(n4916), .CLK(clk), .Q(N3853) );
  DFFPOSX1 \regZ_reg[3][3]  ( .D(n4917), .CLK(clk), .Q(N3856) );
  DFFPOSX1 \regZ_reg[3][2]  ( .D(n4918), .CLK(clk), .Q(N3859) );
  DFFPOSX1 \regZ_reg[3][1]  ( .D(n4919), .CLK(clk), .Q(N3862) );
  DFFPOSX1 \regZ_reg[3][0]  ( .D(n4920), .CLK(clk), .Q(N3865) );
  DFFPOSX1 \regZ_tri_enable_reg[3][0]  ( .D(n4720), .CLK(clk), .Q(N3866) );
  DFFPOSX1 \regZ_tri_enable_reg[3][1]  ( .D(n4719), .CLK(clk), .Q(N3863) );
  DFFPOSX1 \regZ_tri_enable_reg[3][2]  ( .D(n4718), .CLK(clk), .Q(N3860) );
  DFFPOSX1 \regZ_tri_enable_reg[3][3]  ( .D(n4717), .CLK(clk), .Q(N3857) );
  DFFPOSX1 \regZ_tri_enable_reg[3][4]  ( .D(n4716), .CLK(clk), .Q(N3854) );
  DFFPOSX1 \regZ_tri_enable_reg[3][5]  ( .D(n4715), .CLK(clk), .Q(N3851) );
  DFFPOSX1 \regZ_tri_enable_reg[3][6]  ( .D(n4714), .CLK(clk), .Q(N3848) );
  DFFPOSX1 \regZ_tri_enable_reg[3][7]  ( .D(n4713), .CLK(clk), .Q(N3845) );
  DFFPOSX1 \regZ_reg[0][3]  ( .D(n4889), .CLK(clk), .Q(N3784) );
  DFFPOSX1 \regZ_reg[0][2]  ( .D(n4890), .CLK(clk), .Q(N3787) );
  DFFPOSX1 \regZ_reg[0][1]  ( .D(n4891), .CLK(clk), .Q(N3790) );
  DFFPOSX1 \regZ_reg[0][0]  ( .D(n4892), .CLK(clk), .Q(N3793) );
  DFFPOSX1 \regZ_reg[0][7]  ( .D(n4893), .CLK(clk), .Q(N3772) );
  DFFPOSX1 \regZ_reg[0][6]  ( .D(n4894), .CLK(clk), .Q(N3775) );
  DFFPOSX1 \regZ_reg[0][5]  ( .D(n4895), .CLK(clk), .Q(N3778) );
  DFFPOSX1 \regZ_reg[0][4]  ( .D(n4896), .CLK(clk), .Q(N3781) );
  DFFPOSX1 \regZ_tri_enable_reg[0][0]  ( .D(n4696), .CLK(clk), .Q(N3794) );
  DFFPOSX1 \regZ_tri_enable_reg[0][1]  ( .D(n4695), .CLK(clk), .Q(N3791) );
  DFFPOSX1 \regZ_tri_enable_reg[0][2]  ( .D(n4694), .CLK(clk), .Q(N3788) );
  DFFPOSX1 \regZ_tri_enable_reg[0][3]  ( .D(n4693), .CLK(clk), .Q(N3785) );
  DFFPOSX1 \regZ_tri_enable_reg[0][4]  ( .D(n4692), .CLK(clk), .Q(N3782) );
  DFFPOSX1 \regZ_tri_enable_reg[0][5]  ( .D(n4691), .CLK(clk), .Q(N3779) );
  DFFPOSX1 \regZ_tri_enable_reg[0][6]  ( .D(n4690), .CLK(clk), .Q(N3776) );
  DFFPOSX1 \regZ_tri_enable_reg[0][7]  ( .D(n4689), .CLK(clk), .Q(N3773) );
  DFFPOSX1 \Out_bThres_reg[0]  ( .D(n4652), .CLK(clk), .Q(\Out_bThres[0] ) );
  DFFPOSX1 \Out_gradient_reg[7]  ( .D(n4661), .CLK(clk), .Q(N4396) );
  DFFPOSX1 \Out_gradient_reg[6]  ( .D(n4662), .CLK(clk), .Q(N4399) );
  DFFPOSX1 \Out_gradient_reg[5]  ( .D(n4663), .CLK(clk), .Q(N4402) );
  DFFPOSX1 \Out_gradient_reg[4]  ( .D(n4664), .CLK(clk), .Q(N4405) );
  DFFPOSX1 \Out_gradient_reg[3]  ( .D(n4665), .CLK(clk), .Q(N4408) );
  DFFPOSX1 \Out_gradient_reg[2]  ( .D(n4666), .CLK(clk), .Q(N4411) );
  DFFPOSX1 \Out_gradient_reg[1]  ( .D(n4667), .CLK(clk), .Q(N4414) );
  DFFPOSX1 \Out_gradient_reg[0]  ( .D(n4668), .CLK(clk), .Q(N4417) );
  DFFPOSX1 \Out_gradient_tri_enable_reg[7]  ( .D(n4669), .CLK(clk), .Q(N4397)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[6]  ( .D(n4670), .CLK(clk), .Q(N4400)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[5]  ( .D(n4671), .CLK(clk), .Q(N4403)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[4]  ( .D(n4672), .CLK(clk), .Q(N4406)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[3]  ( .D(n4673), .CLK(clk), .Q(N4409)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[2]  ( .D(n4674), .CLK(clk), .Q(N4412)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[1]  ( .D(n4675), .CLK(clk), .Q(N4415)
         );
  DFFPOSX1 \Out_gradient_tri_enable_reg[0]  ( .D(n4676), .CLK(clk), .Q(N4418)
         );
  DFFPOSX1 \Out_direction_reg[7]  ( .D(n4637), .CLK(clk), .Q(N4420) );
  DFFPOSX1 \Out_direction_reg[2]  ( .D(n4647), .CLK(clk), .Q(N4435) );
  DFFPOSX1 \Out_direction_reg[0]  ( .D(n4651), .CLK(clk), .Q(N4441) );
  DFFPOSX1 \Out_direction_tri_enable_reg[0]  ( .D(n4650), .CLK(clk), .Q(N4442)
         );
  DFFPOSX1 \Out_direction_reg[1]  ( .D(n4649), .CLK(clk), .Q(N4438) );
  DFFPOSX1 \Out_direction_tri_enable_reg[1]  ( .D(n4648), .CLK(clk), .Q(N4439)
         );
  DFFPOSX1 \Out_direction_tri_enable_reg[2]  ( .D(n4646), .CLK(clk), .Q(N4436)
         );
  DFFPOSX1 \Out_direction_reg[3]  ( .D(n4645), .CLK(clk), .Q(N4432) );
  DFFPOSX1 \Out_direction_tri_enable_reg[3]  ( .D(n4644), .CLK(clk), .Q(N4433)
         );
  DFFPOSX1 \Out_direction_reg[4]  ( .D(n4643), .CLK(clk), .Q(N4429) );
  DFFPOSX1 \Out_direction_tri_enable_reg[4]  ( .D(n4642), .CLK(clk), .Q(N4430)
         );
  DFFPOSX1 \Out_direction_reg[5]  ( .D(n4641), .CLK(clk), .Q(N4426) );
  DFFPOSX1 \Out_direction_tri_enable_reg[5]  ( .D(n4640), .CLK(clk), .Q(N4427)
         );
  DFFPOSX1 \Out_direction_reg[6]  ( .D(n4639), .CLK(clk), .Q(N4423) );
  DFFPOSX1 \Out_direction_tri_enable_reg[6]  ( .D(n4638), .CLK(clk), .Q(N4424)
         );
  DFFPOSX1 \Out_direction_tri_enable_reg[7]  ( .D(n4636), .CLK(clk), .Q(N4421)
         );
  DFFPOSX1 \Out_gf_reg[7]  ( .D(n3741), .CLK(clk), .Q(Out_gf[7]) );
  DFFPOSX1 \OutData_reg[7]  ( .D(n4620), .CLK(clk), .Q(N4468) );
  DFFPOSX1 \Out_gf_reg[6]  ( .D(n3742), .CLK(clk), .Q(Out_gf[6]) );
  DFFPOSX1 \OutData_reg[6]  ( .D(n4621), .CLK(clk), .Q(N4471) );
  DFFPOSX1 \Out_gf_reg[5]  ( .D(n3743), .CLK(clk), .Q(Out_gf[5]) );
  DFFPOSX1 \OutData_reg[5]  ( .D(n4622), .CLK(clk), .Q(N4474) );
  DFFPOSX1 \Out_gf_reg[4]  ( .D(n3744), .CLK(clk), .Q(Out_gf[4]) );
  DFFPOSX1 \OutData_reg[4]  ( .D(n4623), .CLK(clk), .Q(N4477) );
  DFFPOSX1 \Out_gf_reg[3]  ( .D(n3745), .CLK(clk), .Q(Out_gf[3]) );
  DFFPOSX1 \OutData_reg[3]  ( .D(n4624), .CLK(clk), .Q(N4480) );
  DFFPOSX1 \Out_gf_reg[2]  ( .D(n3746), .CLK(clk), .Q(Out_gf[2]) );
  DFFPOSX1 \OutData_reg[2]  ( .D(n4625), .CLK(clk), .Q(N4483) );
  DFFPOSX1 \Out_gf_reg[1]  ( .D(n3747), .CLK(clk), .Q(Out_gf[1]) );
  DFFPOSX1 \OutData_reg[1]  ( .D(n4626), .CLK(clk), .Q(N4486) );
  DFFPOSX1 \Out_gf_reg[0]  ( .D(n3748), .CLK(clk), .Q(Out_gf[0]) );
  DFFPOSX1 \OutData_reg[0]  ( .D(n4627), .CLK(clk), .Q(N4489) );
  TBUFX1 \dx_tri[0]  ( .A(n7279), .EN(n7278), .Y(dx[0]) );
  TBUFX1 \dy_tri[0]  ( .A(n7280), .EN(n7281), .Y(dy[0]) );
  TBUFX1 \OutData_tri[0]  ( .A(n7737), .EN(n7261), .Y(OutData[0]) );
  TBUFX1 \OutData_tri[1]  ( .A(n7736), .EN(n7260), .Y(OutData[1]) );
  TBUFX1 \OutData_tri[2]  ( .A(n7735), .EN(n7259), .Y(OutData[2]) );
  TBUFX1 \OutData_tri[3]  ( .A(n7734), .EN(n7258), .Y(OutData[3]) );
  TBUFX1 \OutData_tri[4]  ( .A(n7733), .EN(n7257), .Y(OutData[4]) );
  TBUFX1 \OutData_tri[5]  ( .A(n7732), .EN(n7256), .Y(OutData[5]) );
  TBUFX1 \OutData_tri[6]  ( .A(n7731), .EN(n7255), .Y(OutData[6]) );
  TBUFX1 \OutData_tri[7]  ( .A(n7730), .EN(n7254), .Y(OutData[7]) );
  TBUFX1 \fGy_tri[0]  ( .A(n7283), .EN(n7270), .Y(fGy[0]) );
  TBUFX1 \fGy_tri[1]  ( .A(n7284), .EN(n7271), .Y(fGy[1]) );
  TBUFX1 \fGy_tri[2]  ( .A(n7285), .EN(n7272), .Y(fGy[2]) );
  TBUFX1 \fGy_tri[3]  ( .A(n7286), .EN(n7273), .Y(fGy[3]) );
  TBUFX1 \fGy_tri[4]  ( .A(n7287), .EN(n7274), .Y(fGy[4]) );
  TBUFX1 \fGy_tri[5]  ( .A(n7288), .EN(n7275), .Y(fGy[5]) );
  TBUFX1 \fGy_tri[6]  ( .A(n7289), .EN(n7276), .Y(fGy[6]) );
  TBUFX1 \fGy_tri[7]  ( .A(n7290), .EN(n7277), .Y(fGy[7]) );
  TBUFX1 \Out_direction_tri[0]  ( .A(n7716), .EN(n7717), .Y(Out_direction[0])
         );
  TBUFX1 \Out_direction_tri[1]  ( .A(n7718), .EN(n7719), .Y(Out_direction[1])
         );
  TBUFX1 \Out_direction_tri[2]  ( .A(n7715), .EN(n7720), .Y(Out_direction[2])
         );
  TBUFX1 \Out_direction_tri[3]  ( .A(n7721), .EN(n7722), .Y(Out_direction[3])
         );
  TBUFX1 \Out_direction_tri[4]  ( .A(n7723), .EN(n7724), .Y(Out_direction[4])
         );
  TBUFX1 \Out_direction_tri[5]  ( .A(n7725), .EN(n7726), .Y(Out_direction[5])
         );
  TBUFX1 \Out_direction_tri[6]  ( .A(n7727), .EN(n7728), .Y(Out_direction[6])
         );
  TBUFX1 \Out_direction_tri[7]  ( .A(n7714), .EN(n7729), .Y(Out_direction[7])
         );
  TBUFX1 \Out_gradient_tri[0]  ( .A(n7705), .EN(n7713), .Y(Out_gradient[0]) );
  TBUFX1 \Out_gradient_tri[1]  ( .A(n7704), .EN(n7712), .Y(Out_gradient[1]) );
  TBUFX1 \Out_gradient_tri[2]  ( .A(n7703), .EN(n7711), .Y(Out_gradient[2]) );
  TBUFX1 \Out_gradient_tri[3]  ( .A(n7702), .EN(n7710), .Y(Out_gradient[3]) );
  TBUFX1 \Out_gradient_tri[4]  ( .A(n7701), .EN(n7709), .Y(Out_gradient[4]) );
  TBUFX1 \Out_gradient_tri[5]  ( .A(n7700), .EN(n7708), .Y(Out_gradient[5]) );
  TBUFX1 \Out_gradient_tri[6]  ( .A(n7699), .EN(n7707), .Y(Out_gradient[6]) );
  TBUFX1 \Out_gradient_tri[7]  ( .A(n7698), .EN(n7706), .Y(Out_gradient[7]) );
  TBUFX1 \fGx_tri[0]  ( .A(n7282), .EN(n7262), .Y(fGx[0]) );
  TBUFX1 \fGx_tri[1]  ( .A(n7291), .EN(n7263), .Y(fGx[1]) );
  TBUFX1 \fGx_tri[2]  ( .A(n7292), .EN(n7264), .Y(fGx[2]) );
  TBUFX1 \fGx_tri[3]  ( .A(n7293), .EN(n7265), .Y(fGx[3]) );
  TBUFX1 \fGx_tri[4]  ( .A(n7294), .EN(n7266), .Y(fGx[4]) );
  TBUFX1 \fGx_tri[5]  ( .A(n7295), .EN(n7267), .Y(fGx[5]) );
  TBUFX1 \fGx_tri[6]  ( .A(n7296), .EN(n7268), .Y(fGx[6]) );
  TBUFX1 \fGx_tri[7]  ( .A(n7297), .EN(n7269), .Y(fGx[7]) );
  TBUFX1 \regZ_tri[24][0]  ( .A(n7529), .EN(n7530), .Y(\regZ[24][0] ) );
  TBUFX1 \regZ_tri[24][1]  ( .A(n7528), .EN(n7531), .Y(\regZ[24][1] ) );
  TBUFX1 \regZ_tri[24][2]  ( .A(n7527), .EN(n7532), .Y(\regZ[24][2] ) );
  TBUFX1 \regZ_tri[24][3]  ( .A(n7526), .EN(n7533), .Y(\regZ[24][3] ) );
  TBUFX1 \regZ_tri[24][4]  ( .A(n7525), .EN(n7534), .Y(\regZ[24][4] ) );
  TBUFX1 \regZ_tri[24][5]  ( .A(n7524), .EN(n7535), .Y(\regZ[24][5] ) );
  TBUFX1 \regZ_tri[24][6]  ( .A(n7523), .EN(n7536), .Y(\regZ[24][6] ) );
  TBUFX1 \regZ_tri[24][7]  ( .A(n7522), .EN(n7537), .Y(\regZ[24][7] ) );
  TBUFX1 \regZ_tri[23][0]  ( .A(n7506), .EN(n7521), .Y(\regZ[23][0] ) );
  TBUFX1 \regZ_tri[23][1]  ( .A(n7507), .EN(n7520), .Y(\regZ[23][1] ) );
  TBUFX1 \regZ_tri[23][2]  ( .A(n7508), .EN(n7519), .Y(\regZ[23][2] ) );
  TBUFX1 \regZ_tri[23][3]  ( .A(n7509), .EN(n7518), .Y(\regZ[23][3] ) );
  TBUFX1 \regZ_tri[23][4]  ( .A(n7510), .EN(n7517), .Y(\regZ[23][4] ) );
  TBUFX1 \regZ_tri[23][5]  ( .A(n7511), .EN(n7516), .Y(\regZ[23][5] ) );
  TBUFX1 \regZ_tri[23][6]  ( .A(n7512), .EN(n7515), .Y(\regZ[23][6] ) );
  TBUFX1 \regZ_tri[23][7]  ( .A(n7513), .EN(n7514), .Y(\regZ[23][7] ) );
  TBUFX1 \regZ_tri[22][0]  ( .A(n7490), .EN(n7505), .Y(\regZ[22][0] ) );
  TBUFX1 \regZ_tri[22][1]  ( .A(n7491), .EN(n7504), .Y(\regZ[22][1] ) );
  TBUFX1 \regZ_tri[22][2]  ( .A(n7492), .EN(n7503), .Y(\regZ[22][2] ) );
  TBUFX1 \regZ_tri[22][3]  ( .A(n7493), .EN(n7502), .Y(\regZ[22][3] ) );
  TBUFX1 \regZ_tri[22][4]  ( .A(n7494), .EN(n7501), .Y(\regZ[22][4] ) );
  TBUFX1 \regZ_tri[22][5]  ( .A(n7495), .EN(n7500), .Y(\regZ[22][5] ) );
  TBUFX1 \regZ_tri[22][6]  ( .A(n7496), .EN(n7499), .Y(\regZ[22][6] ) );
  TBUFX1 \regZ_tri[22][7]  ( .A(n7497), .EN(n7498), .Y(\regZ[22][7] ) );
  TBUFX1 \regZ_tri[21][0]  ( .A(n7442), .EN(n7457), .Y(\regZ[21][0] ) );
  TBUFX1 \regZ_tri[21][1]  ( .A(n7443), .EN(n7456), .Y(\regZ[21][1] ) );
  TBUFX1 \regZ_tri[21][2]  ( .A(n7444), .EN(n7455), .Y(\regZ[21][2] ) );
  TBUFX1 \regZ_tri[21][3]  ( .A(n7445), .EN(n7454), .Y(\regZ[21][3] ) );
  TBUFX1 \regZ_tri[21][4]  ( .A(n7446), .EN(n7453), .Y(\regZ[21][4] ) );
  TBUFX1 \regZ_tri[21][5]  ( .A(n7447), .EN(n7452), .Y(\regZ[21][5] ) );
  TBUFX1 \regZ_tri[21][6]  ( .A(n7448), .EN(n7451), .Y(\regZ[21][6] ) );
  TBUFX1 \regZ_tri[21][7]  ( .A(n7449), .EN(n7450), .Y(\regZ[21][7] ) );
  TBUFX1 \regZ_tri[20][0]  ( .A(n7426), .EN(n7441), .Y(\regZ[20][0] ) );
  TBUFX1 \regZ_tri[20][1]  ( .A(n7427), .EN(n7440), .Y(\regZ[20][1] ) );
  TBUFX1 \regZ_tri[20][2]  ( .A(n7428), .EN(n7439), .Y(\regZ[20][2] ) );
  TBUFX1 \regZ_tri[20][3]  ( .A(n7429), .EN(n7438), .Y(\regZ[20][3] ) );
  TBUFX1 \regZ_tri[20][4]  ( .A(n7430), .EN(n7437), .Y(\regZ[20][4] ) );
  TBUFX1 \regZ_tri[20][5]  ( .A(n7431), .EN(n7436), .Y(\regZ[20][5] ) );
  TBUFX1 \regZ_tri[20][6]  ( .A(n7432), .EN(n7435), .Y(\regZ[20][6] ) );
  TBUFX1 \regZ_tri[20][7]  ( .A(n7433), .EN(n7434), .Y(\regZ[20][7] ) );
  TBUFX1 \regZ_tri[19][0]  ( .A(n7378), .EN(n7393), .Y(\regZ[19][0] ) );
  TBUFX1 \regZ_tri[19][1]  ( .A(n7379), .EN(n7392), .Y(\regZ[19][1] ) );
  TBUFX1 \regZ_tri[19][2]  ( .A(n7380), .EN(n7391), .Y(\regZ[19][2] ) );
  TBUFX1 \regZ_tri[19][3]  ( .A(n7381), .EN(n7390), .Y(\regZ[19][3] ) );
  TBUFX1 \regZ_tri[19][4]  ( .A(n7382), .EN(n7389), .Y(\regZ[19][4] ) );
  TBUFX1 \regZ_tri[19][5]  ( .A(n7383), .EN(n7388), .Y(\regZ[19][5] ) );
  TBUFX1 \regZ_tri[19][6]  ( .A(n7384), .EN(n7387), .Y(\regZ[19][6] ) );
  TBUFX1 \regZ_tri[19][7]  ( .A(n7385), .EN(n7386), .Y(\regZ[19][7] ) );
  TBUFX1 \regZ_tri[18][0]  ( .A(n7362), .EN(n7377), .Y(\regZ[18][0] ) );
  TBUFX1 \regZ_tri[18][1]  ( .A(n7363), .EN(n7376), .Y(\regZ[18][1] ) );
  TBUFX1 \regZ_tri[18][2]  ( .A(n7364), .EN(n7375), .Y(\regZ[18][2] ) );
  TBUFX1 \regZ_tri[18][3]  ( .A(n7365), .EN(n7374), .Y(\regZ[18][3] ) );
  TBUFX1 \regZ_tri[18][4]  ( .A(n7366), .EN(n7373), .Y(\regZ[18][4] ) );
  TBUFX1 \regZ_tri[18][5]  ( .A(n7367), .EN(n7372), .Y(\regZ[18][5] ) );
  TBUFX1 \regZ_tri[18][6]  ( .A(n7368), .EN(n7371), .Y(\regZ[18][6] ) );
  TBUFX1 \regZ_tri[18][7]  ( .A(n7369), .EN(n7370), .Y(\regZ[18][7] ) );
  TBUFX1 \regZ_tri[17][0]  ( .A(n7545), .EN(n7546), .Y(\regZ[17][0] ) );
  TBUFX1 \regZ_tri[17][1]  ( .A(n7544), .EN(n7547), .Y(\regZ[17][1] ) );
  TBUFX1 \regZ_tri[17][2]  ( .A(n7543), .EN(n7548), .Y(\regZ[17][2] ) );
  TBUFX1 \regZ_tri[17][3]  ( .A(n7542), .EN(n7549), .Y(\regZ[17][3] ) );
  TBUFX1 \regZ_tri[17][4]  ( .A(n7541), .EN(n7550), .Y(\regZ[17][4] ) );
  TBUFX1 \regZ_tri[17][5]  ( .A(n7540), .EN(n7551), .Y(\regZ[17][5] ) );
  TBUFX1 \regZ_tri[17][6]  ( .A(n7539), .EN(n7552), .Y(\regZ[17][6] ) );
  TBUFX1 \regZ_tri[17][7]  ( .A(n7538), .EN(n7553), .Y(\regZ[17][7] ) );
  TBUFX1 \regZ_tri[16][0]  ( .A(n7561), .EN(n7562), .Y(\regZ[16][0] ) );
  TBUFX1 \regZ_tri[16][1]  ( .A(n7560), .EN(n7563), .Y(\regZ[16][1] ) );
  TBUFX1 \regZ_tri[16][2]  ( .A(n7559), .EN(n7564), .Y(\regZ[16][2] ) );
  TBUFX1 \regZ_tri[16][3]  ( .A(n7558), .EN(n7565), .Y(\regZ[16][3] ) );
  TBUFX1 \regZ_tri[16][4]  ( .A(n7557), .EN(n7566), .Y(\regZ[16][4] ) );
  TBUFX1 \regZ_tri[16][5]  ( .A(n7556), .EN(n7567), .Y(\regZ[16][5] ) );
  TBUFX1 \regZ_tri[16][6]  ( .A(n7555), .EN(n7568), .Y(\regZ[16][6] ) );
  TBUFX1 \regZ_tri[16][7]  ( .A(n7554), .EN(n7569), .Y(\regZ[16][7] ) );
  TBUFX1 \regZ_tri[15][0]  ( .A(n7474), .EN(n7489), .Y(\regZ[15][0] ) );
  TBUFX1 \regZ_tri[15][1]  ( .A(n7475), .EN(n7488), .Y(\regZ[15][1] ) );
  TBUFX1 \regZ_tri[15][2]  ( .A(n7476), .EN(n7487), .Y(\regZ[15][2] ) );
  TBUFX1 \regZ_tri[15][3]  ( .A(n7477), .EN(n7486), .Y(\regZ[15][3] ) );
  TBUFX1 \regZ_tri[15][4]  ( .A(n7478), .EN(n7485), .Y(\regZ[15][4] ) );
  TBUFX1 \regZ_tri[15][5]  ( .A(n7479), .EN(n7484), .Y(\regZ[15][5] ) );
  TBUFX1 \regZ_tri[15][6]  ( .A(n7480), .EN(n7483), .Y(\regZ[15][6] ) );
  TBUFX1 \regZ_tri[15][7]  ( .A(n7481), .EN(n7482), .Y(\regZ[15][7] ) );
  TBUFX1 \regZ_tri[14][0]  ( .A(n7458), .EN(n7473), .Y(\regZ[14][0] ) );
  TBUFX1 \regZ_tri[14][1]  ( .A(n7459), .EN(n7472), .Y(\regZ[14][1] ) );
  TBUFX1 \regZ_tri[14][2]  ( .A(n7460), .EN(n7471), .Y(\regZ[14][2] ) );
  TBUFX1 \regZ_tri[14][3]  ( .A(n7461), .EN(n7470), .Y(\regZ[14][3] ) );
  TBUFX1 \regZ_tri[14][4]  ( .A(n7462), .EN(n7469), .Y(\regZ[14][4] ) );
  TBUFX1 \regZ_tri[14][5]  ( .A(n7463), .EN(n7468), .Y(\regZ[14][5] ) );
  TBUFX1 \regZ_tri[14][6]  ( .A(n7464), .EN(n7467), .Y(\regZ[14][6] ) );
  TBUFX1 \regZ_tri[14][7]  ( .A(n7465), .EN(n7466), .Y(\regZ[14][7] ) );
  TBUFX1 \regZ_tri[13][0]  ( .A(n7410), .EN(n7425), .Y(\regZ[13][0] ) );
  TBUFX1 \regZ_tri[13][1]  ( .A(n7411), .EN(n7424), .Y(\regZ[13][1] ) );
  TBUFX1 \regZ_tri[13][2]  ( .A(n7412), .EN(n7423), .Y(\regZ[13][2] ) );
  TBUFX1 \regZ_tri[13][3]  ( .A(n7413), .EN(n7422), .Y(\regZ[13][3] ) );
  TBUFX1 \regZ_tri[13][4]  ( .A(n7414), .EN(n7421), .Y(\regZ[13][4] ) );
  TBUFX1 \regZ_tri[13][5]  ( .A(n7415), .EN(n7420), .Y(\regZ[13][5] ) );
  TBUFX1 \regZ_tri[13][6]  ( .A(n7416), .EN(n7419), .Y(\regZ[13][6] ) );
  TBUFX1 \regZ_tri[13][7]  ( .A(n7417), .EN(n7418), .Y(\regZ[13][7] ) );
  TBUFX1 \regZ_tri[12][0]  ( .A(n7394), .EN(n7402), .Y(\regZ[12][0] ) );
  TBUFX1 \regZ_tri[12][1]  ( .A(n7401), .EN(n7403), .Y(\regZ[12][1] ) );
  TBUFX1 \regZ_tri[12][2]  ( .A(n7400), .EN(n7404), .Y(\regZ[12][2] ) );
  TBUFX1 \regZ_tri[12][3]  ( .A(n7399), .EN(n7405), .Y(\regZ[12][3] ) );
  TBUFX1 \regZ_tri[12][4]  ( .A(n7398), .EN(n7406), .Y(\regZ[12][4] ) );
  TBUFX1 \regZ_tri[12][5]  ( .A(n7397), .EN(n7407), .Y(\regZ[12][5] ) );
  TBUFX1 \regZ_tri[12][6]  ( .A(n7396), .EN(n7408), .Y(\regZ[12][6] ) );
  TBUFX1 \regZ_tri[12][7]  ( .A(n7395), .EN(n7409), .Y(\regZ[12][7] ) );
  TBUFX1 \regZ_tri[11][0]  ( .A(n7346), .EN(n7361), .Y(\regZ[11][0] ) );
  TBUFX1 \regZ_tri[11][1]  ( .A(n7347), .EN(n7360), .Y(\regZ[11][1] ) );
  TBUFX1 \regZ_tri[11][2]  ( .A(n7348), .EN(n7359), .Y(\regZ[11][2] ) );
  TBUFX1 \regZ_tri[11][3]  ( .A(n7349), .EN(n7358), .Y(\regZ[11][3] ) );
  TBUFX1 \regZ_tri[11][4]  ( .A(n7350), .EN(n7357), .Y(\regZ[11][4] ) );
  TBUFX1 \regZ_tri[11][5]  ( .A(n7351), .EN(n7356), .Y(\regZ[11][5] ) );
  TBUFX1 \regZ_tri[11][6]  ( .A(n7352), .EN(n7355), .Y(\regZ[11][6] ) );
  TBUFX1 \regZ_tri[11][7]  ( .A(n7353), .EN(n7354), .Y(\regZ[11][7] ) );
  TBUFX1 \regZ_tri[10][0]  ( .A(n7330), .EN(n7345), .Y(\regZ[10][0] ) );
  TBUFX1 \regZ_tri[10][1]  ( .A(n7331), .EN(n7344), .Y(\regZ[10][1] ) );
  TBUFX1 \regZ_tri[10][2]  ( .A(n7332), .EN(n7343), .Y(\regZ[10][2] ) );
  TBUFX1 \regZ_tri[10][3]  ( .A(n7333), .EN(n7342), .Y(\regZ[10][3] ) );
  TBUFX1 \regZ_tri[10][4]  ( .A(n7334), .EN(n7341), .Y(\regZ[10][4] ) );
  TBUFX1 \regZ_tri[10][5]  ( .A(n7335), .EN(n7340), .Y(\regZ[10][5] ) );
  TBUFX1 \regZ_tri[10][6]  ( .A(n7336), .EN(n7339), .Y(\regZ[10][6] ) );
  TBUFX1 \regZ_tri[10][7]  ( .A(n7337), .EN(n7338), .Y(\regZ[10][7] ) );
  TBUFX1 \regZ_tri[9][0]  ( .A(n7577), .EN(n7578), .Y(\regZ[9][0] ) );
  TBUFX1 \regZ_tri[9][1]  ( .A(n7576), .EN(n7579), .Y(\regZ[9][1] ) );
  TBUFX1 \regZ_tri[9][2]  ( .A(n7575), .EN(n7580), .Y(\regZ[9][2] ) );
  TBUFX1 \regZ_tri[9][3]  ( .A(n7574), .EN(n7581), .Y(\regZ[9][3] ) );
  TBUFX1 \regZ_tri[9][4]  ( .A(n7573), .EN(n7582), .Y(\regZ[9][4] ) );
  TBUFX1 \regZ_tri[9][5]  ( .A(n7572), .EN(n7583), .Y(\regZ[9][5] ) );
  TBUFX1 \regZ_tri[9][6]  ( .A(n7571), .EN(n7584), .Y(\regZ[9][6] ) );
  TBUFX1 \regZ_tri[9][7]  ( .A(n7570), .EN(n7585), .Y(\regZ[9][7] ) );
  TBUFX1 \regZ_tri[8][0]  ( .A(n7593), .EN(n7594), .Y(\regZ[8][0] ) );
  TBUFX1 \regZ_tri[8][1]  ( .A(n7592), .EN(n7595), .Y(\regZ[8][1] ) );
  TBUFX1 \regZ_tri[8][2]  ( .A(n7591), .EN(n7596), .Y(\regZ[8][2] ) );
  TBUFX1 \regZ_tri[8][3]  ( .A(n7590), .EN(n7597), .Y(\regZ[8][3] ) );
  TBUFX1 \regZ_tri[8][4]  ( .A(n7589), .EN(n7598), .Y(\regZ[8][4] ) );
  TBUFX1 \regZ_tri[8][5]  ( .A(n7588), .EN(n7599), .Y(\regZ[8][5] ) );
  TBUFX1 \regZ_tri[8][6]  ( .A(n7587), .EN(n7600), .Y(\regZ[8][6] ) );
  TBUFX1 \regZ_tri[8][7]  ( .A(n7586), .EN(n7601), .Y(\regZ[8][7] ) );
  TBUFX1 \regZ_tri[7][0]  ( .A(n7609), .EN(n7610), .Y(\regZ[7][0] ) );
  TBUFX1 \regZ_tri[7][1]  ( .A(n7608), .EN(n7611), .Y(\regZ[7][1] ) );
  TBUFX1 \regZ_tri[7][2]  ( .A(n7607), .EN(n7612), .Y(\regZ[7][2] ) );
  TBUFX1 \regZ_tri[7][3]  ( .A(n7606), .EN(n7613), .Y(\regZ[7][3] ) );
  TBUFX1 \regZ_tri[7][4]  ( .A(n7605), .EN(n7614), .Y(\regZ[7][4] ) );
  TBUFX1 \regZ_tri[7][5]  ( .A(n7604), .EN(n7615), .Y(\regZ[7][5] ) );
  TBUFX1 \regZ_tri[7][6]  ( .A(n7603), .EN(n7616), .Y(\regZ[7][6] ) );
  TBUFX1 \regZ_tri[7][7]  ( .A(n7602), .EN(n7617), .Y(\regZ[7][7] ) );
  TBUFX1 \regZ_tri[6][0]  ( .A(n7625), .EN(n7626), .Y(\regZ[6][0] ) );
  TBUFX1 \regZ_tri[6][1]  ( .A(n7624), .EN(n7627), .Y(\regZ[6][1] ) );
  TBUFX1 \regZ_tri[6][2]  ( .A(n7623), .EN(n7628), .Y(\regZ[6][2] ) );
  TBUFX1 \regZ_tri[6][3]  ( .A(n7622), .EN(n7629), .Y(\regZ[6][3] ) );
  TBUFX1 \regZ_tri[6][4]  ( .A(n7621), .EN(n7630), .Y(\regZ[6][4] ) );
  TBUFX1 \regZ_tri[6][5]  ( .A(n7620), .EN(n7631), .Y(\regZ[6][5] ) );
  TBUFX1 \regZ_tri[6][6]  ( .A(n7619), .EN(n7632), .Y(\regZ[6][6] ) );
  TBUFX1 \regZ_tri[6][7]  ( .A(n7618), .EN(n7633), .Y(\regZ[6][7] ) );
  TBUFX1 \regZ_tri[5][0]  ( .A(n7641), .EN(n7642), .Y(\regZ[5][0] ) );
  TBUFX1 \regZ_tri[5][1]  ( .A(n7640), .EN(n7643), .Y(\regZ[5][1] ) );
  TBUFX1 \regZ_tri[5][2]  ( .A(n7639), .EN(n7644), .Y(\regZ[5][2] ) );
  TBUFX1 \regZ_tri[5][3]  ( .A(n7638), .EN(n7645), .Y(\regZ[5][3] ) );
  TBUFX1 \regZ_tri[5][4]  ( .A(n7637), .EN(n7646), .Y(\regZ[5][4] ) );
  TBUFX1 \regZ_tri[5][5]  ( .A(n7636), .EN(n7647), .Y(\regZ[5][5] ) );
  TBUFX1 \regZ_tri[5][6]  ( .A(n7635), .EN(n7648), .Y(\regZ[5][6] ) );
  TBUFX1 \regZ_tri[5][7]  ( .A(n7634), .EN(n7649), .Y(\regZ[5][7] ) );
  TBUFX1 \regZ_tri[4][0]  ( .A(n7657), .EN(n7658), .Y(\regZ[4][0] ) );
  TBUFX1 \regZ_tri[4][1]  ( .A(n7656), .EN(n7659), .Y(\regZ[4][1] ) );
  TBUFX1 \regZ_tri[4][2]  ( .A(n7655), .EN(n7660), .Y(\regZ[4][2] ) );
  TBUFX1 \regZ_tri[4][3]  ( .A(n7654), .EN(n7661), .Y(\regZ[4][3] ) );
  TBUFX1 \regZ_tri[4][4]  ( .A(n7653), .EN(n7662), .Y(\regZ[4][4] ) );
  TBUFX1 \regZ_tri[4][5]  ( .A(n7652), .EN(n7663), .Y(\regZ[4][5] ) );
  TBUFX1 \regZ_tri[4][6]  ( .A(n7651), .EN(n7664), .Y(\regZ[4][6] ) );
  TBUFX1 \regZ_tri[4][7]  ( .A(n7650), .EN(n7665), .Y(\regZ[4][7] ) );
  TBUFX1 \regZ_tri[3][0]  ( .A(n7673), .EN(n7674), .Y(\regZ[3][0] ) );
  TBUFX1 \regZ_tri[3][1]  ( .A(n7672), .EN(n7675), .Y(\regZ[3][1] ) );
  TBUFX1 \regZ_tri[3][2]  ( .A(n7671), .EN(n7676), .Y(\regZ[3][2] ) );
  TBUFX1 \regZ_tri[3][3]  ( .A(n7670), .EN(n7677), .Y(\regZ[3][3] ) );
  TBUFX1 \regZ_tri[3][4]  ( .A(n7669), .EN(n7678), .Y(\regZ[3][4] ) );
  TBUFX1 \regZ_tri[3][5]  ( .A(n7668), .EN(n7679), .Y(\regZ[3][5] ) );
  TBUFX1 \regZ_tri[3][6]  ( .A(n7667), .EN(n7680), .Y(\regZ[3][6] ) );
  TBUFX1 \regZ_tri[3][7]  ( .A(n7666), .EN(n7681), .Y(\regZ[3][7] ) );
  TBUFX1 \regZ_tri[2][0]  ( .A(n7321), .EN(n7322), .Y(\regZ[2][0] ) );
  TBUFX1 \regZ_tri[2][1]  ( .A(n7320), .EN(n7323), .Y(\regZ[2][1] ) );
  TBUFX1 \regZ_tri[2][2]  ( .A(n7319), .EN(n7324), .Y(\regZ[2][2] ) );
  TBUFX1 \regZ_tri[2][3]  ( .A(n7318), .EN(n7325), .Y(\regZ[2][3] ) );
  TBUFX1 \regZ_tri[2][4]  ( .A(n7317), .EN(n7326), .Y(\regZ[2][4] ) );
  TBUFX1 \regZ_tri[2][5]  ( .A(n7316), .EN(n7327), .Y(\regZ[2][5] ) );
  TBUFX1 \regZ_tri[2][6]  ( .A(n7315), .EN(n7328), .Y(\regZ[2][6] ) );
  TBUFX1 \regZ_tri[2][7]  ( .A(n7314), .EN(n7329), .Y(\regZ[2][7] ) );
  TBUFX1 \regZ_tri[1][0]  ( .A(n7305), .EN(n7306), .Y(\regZ[1][0] ) );
  TBUFX1 \regZ_tri[1][1]  ( .A(n7304), .EN(n7307), .Y(\regZ[1][1] ) );
  TBUFX1 \regZ_tri[1][2]  ( .A(n7303), .EN(n7308), .Y(\regZ[1][2] ) );
  TBUFX1 \regZ_tri[1][3]  ( .A(n7302), .EN(n7309), .Y(\regZ[1][3] ) );
  TBUFX1 \regZ_tri[1][4]  ( .A(n7301), .EN(n7310), .Y(\regZ[1][4] ) );
  TBUFX1 \regZ_tri[1][5]  ( .A(n7300), .EN(n7311), .Y(\regZ[1][5] ) );
  TBUFX1 \regZ_tri[1][6]  ( .A(n7299), .EN(n7312), .Y(\regZ[1][6] ) );
  TBUFX1 \regZ_tri[1][7]  ( .A(n7298), .EN(n7313), .Y(\regZ[1][7] ) );
  TBUFX1 \regZ_tri[0][0]  ( .A(n7685), .EN(n7690), .Y(\regZ[0][0] ) );
  TBUFX1 \regZ_tri[0][1]  ( .A(n7684), .EN(n7691), .Y(\regZ[0][1] ) );
  TBUFX1 \regZ_tri[0][2]  ( .A(n7683), .EN(n7692), .Y(\regZ[0][2] ) );
  TBUFX1 \regZ_tri[0][3]  ( .A(n7682), .EN(n7693), .Y(\regZ[0][3] ) );
  TBUFX1 \regZ_tri[0][4]  ( .A(n7689), .EN(n7694), .Y(\regZ[0][4] ) );
  TBUFX1 \regZ_tri[0][5]  ( .A(n7688), .EN(n7695), .Y(\regZ[0][5] ) );
  TBUFX1 \regZ_tri[0][6]  ( .A(n7687), .EN(n7696), .Y(\regZ[0][6] ) );
  TBUFX1 \regZ_tri[0][7]  ( .A(n7686), .EN(n7697), .Y(\regZ[0][7] ) );
  CannyEdge_DW01_addsub_1 add_0_root_add_205_8 ( .A({N2416, N2415, N2414, 
        N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, 
        N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, 
        N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385}), .B({
        N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, 
        N2470, N2469, N2468, N2467, N2466, N2465, N2464, N1912, N1911, N1910, 
        N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, 
        N1899, N1898}), .CI(1'b0), .ADD_SUB(1'b0), .SUM({N2544, N2543, N2542, 
        N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, 
        N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, 
        N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513}) );
  CannyEdge_DW01_addsub_3 add_0_root_add_160_24 ( .A({N2002, N2001, N2000, 
        N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, 
        N1989, N1988}), .B({N2032, N2031, N2030, N2029, N2028, N2027, N2026, 
        N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N2055, N2054, N2053, N2052, N2051, N2050, N2049, 
        N2048, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  CannyEdge_DW01_addsub_4 add_1_root_add_160_24 ( .A({N1942, N1941, N1940, 
        N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, 
        N1929, N1928}), .B({N1972, N1971, N1970, N1969, N1968, N1967, N1966, 
        N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N2032, N2031, N2030, N2029, N2028, N2027, N2026, 
        N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018}) );
  CannyEdge_DW01_add_0 add_3_root_add_160_24 ( .A({N1822, N1821, N1820, N1819, 
        N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, 
        1'b0}), .B({N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, 
        N1844, N1843, N1842, N1841, N1840, N1839, N1838}), .CI(1'b0), .SUM({
        N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, 
        N1962, N1961, N1960, N1959, N1958}) );
  CannyEdge_DW01_add_1 add_7_root_add_160_24 ( .A({N1582, N1581, N1580, N1579, 
        N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, 
        N1568}), .B({N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, 
        N1604, N1603, N1602, N1601, N1600, N1599, N1598}), .CI(1'b0), .SUM({
        N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, 
        N1842, N1841, N1840, N1839, N1838}) );
  CannyEdge_DW01_add_2 add_15_root_add_160_24 ( .A({1'b0, N1806, N1805, N1804, 
        N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, 
        N1793}), .B({1'b0, N1836, N1835, N1834, N1833, N1832, N1831, N1830, 
        N1829, N1828, N1827, N1826, N1825, N1824, 1'b0}), .CI(1'b0), .SUM({
        N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, 
        N1602, N1601, N1600, N1599, N1598}) );
  CannyEdge_DW01_add_4 add_8_root_add_160_24 ( .A({N1522, N1521, N1520, N1519, 
        N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, 
        1'b0}), .B({N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, 
        N1544, N1543, N1542, N1541, N1540, N1539, 1'b0}), .CI(1'b0), .SUM({
        N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, 
        N1812, N1811, N1810, N1809, SYNOPSYS_UNCONNECTED__7}) );
  CannyEdge_DW01_add_7 add_4_root_add_160_24 ( .A({N1762, N1761, N1760, N1759, 
        N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, 
        N1748}), .B({N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, 
        N1784, N1783, N1782, N1781, N1780, N1779, N1778}), .CI(1'b0), .SUM({
        N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, 
        N1932, N1931, N1930, N1929, N1928}) );
  CannyEdge_DW01_add_8 add_9_root_add_160_24 ( .A({N1462, N1461, N1460, N1459, 
        N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, 
        N1448}), .B({N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, 
        N1484, N1483, N1482, N1481, N1480, N1479, N1478}), .CI(1'b0), .SUM({
        N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, 
        N1782, N1781, N1780, N1779, N1778}) );
  CannyEdge_DW01_add_9 add_19_root_add_160_24 ( .A({1'b0, N1566, N1565, N1564, 
        N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, 
        N1553}), .B({1'b0, N1596, N1595, N1594, N1593, N1592, N1591, N1590, 
        N1589, N1588, N1587, N1586, N1585, N1584, N1583}), .CI(1'b0), .SUM({
        N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, 
        N1482, N1481, N1480, N1479, N1478}) );
  CannyEdge_DW01_add_10 add_10_root_add_160_24 ( .A({N1402, N1401, N1400, 
        N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, 
        N1389, N1388}), .B({N2186, N2185, N2184, N2183, N2182, N2181, N2180, 
        N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172}), .CI(1'b0), 
        .SUM({N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, 
        N1753, N1752, N1751, N1750, N1749, N1748}) );
  CannyEdge_DW01_add_11 add_2_root_add_160_24 ( .A({N1882, N1881, N1880, N1879, 
        N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, 
        N1868}), .B({N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, 
        N1904, N1903, N1902, N1901, N1900, N1899, N1898}), .CI(1'b0), .SUM({
        N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, 
        N1992, N1991, N1990, N1989, N1988}) );
  CannyEdge_DW01_add_12 r1417 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U76/Z_14 , \U3/U76/Z_13 , \U3/U76/Z_12 , \U3/U76/Z_11 , 
        \U3/U76/Z_10 , n7206, n7207, n7208, n7233, n7234, n7235, n7236, n7237, 
        n7238, n7239}), .B({\U3/U77/Z_31 , \U3/U77/Z_30 , \U3/U77/Z_29 , 
        \U3/U77/Z_28 , \U3/U77/Z_27 , \U3/U77/Z_26 , \U3/U77/Z_25 , 
        \U3/U77/Z_24 , \U3/U77/Z_23 , \U3/U77/Z_22 , \U3/U77/Z_21 , 
        \U3/U77/Z_20 , \U3/U77/Z_19 , \U3/U77/Z_18 , \U3/U77/Z_17 , 
        \U3/U77/Z_16 , \U3/U77/Z_15 , N1732, N1731, N1730, N1729, N1728, N1727, 
        N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718}), .CI(
        1'b0), .SUM({N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, 
        N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N1912, 
        N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, 
        N1901, N1900, N1899, N1898}) );
  CannyEdge_DW01_add_13 add_4_root_add_205_8 ( .A({1'b0, 1'b0, \regX[0][7] , 
        \regX[0][6] , \regX[0][5] , \regX[0][4] , \regX[0][3] , \regX[0][2] , 
        \regX[0][1] , \regX[0][0] }), .B({1'b0, \regX[1][7] , \regX[1][6] , 
        \regX[1][5] , \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] , 
        \regX[1][0] , 1'b0}), .CI(1'b0), .SUM({N2341, N2340, N2339, N2338, 
        N2337, N2336, N2335, N2334, N2333, N2332}) );
  CannyEdge_DW01_add_14 r1263 ( .A({\U3/U74/Z_31 , \U3/U74/Z_30 , 
        \U3/U74/Z_29 , \U3/U74/Z_28 , \U3/U74/Z_27 , \U3/U74/Z_26 , 
        \U3/U74/Z_25 , \U3/U74/Z_24 , \U3/U74/Z_23 , \U3/U74/Z_22 , 
        \U3/U74/Z_21 , \U3/U74/Z_20 , \U3/U74/Z_19 , \U3/U74/Z_18 , 
        \U3/U74/Z_17 , \U3/U74/Z_16 , \U3/U74/Z_15 , N2250, N2249, N2248, 
        N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, 
        N2237, N2236}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \U3/U75/Z_14 , 
        \U3/U75/Z_13 , \U3/U75/Z_12 , \U3/U75/Z_11 , \U3/U75/Z_10 , 
        \U3/U75/Z_9 , \U3/U75/Z_8 , \U3/U75/Z_7 , \U3/U75/Z_6 , \U3/U75/Z_5 , 
        \U3/U75/Z_4 , \U3/U75/Z_3 , \U3/U75/Z_2 , \U3/U75/Z_1 , \U3/U75/Z_0 }), 
        .CI(1'b0), .SUM({\U3/U77/DATA2_31 , \U3/U77/DATA2_30 , 
        \U3/U77/DATA2_29 , \U3/U77/DATA2_28 , \U3/U77/DATA2_27 , 
        \U3/U77/DATA2_26 , \U3/U77/DATA2_25 , \U3/U77/DATA2_24 , 
        \U3/U77/DATA2_23 , \U3/U77/DATA2_22 , \U3/U77/DATA2_21 , 
        \U3/U77/DATA2_20 , \U3/U77/DATA2_19 , \U3/U77/DATA2_18 , 
        \U3/U77/DATA2_17 , \U3/U77/DATA2_16 , \U3/U77/DATA2_15 , N1732, N1731, 
        N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, 
        N1720, N1719, N1718}) );
  CannyEdge_DW01_add_15 r1259 ( .A({\U3/U72/Z_31 , \U3/U72/Z_30 , 
        \U3/U72/Z_29 , \U3/U72/Z_28 , \U3/U72/Z_27 , \U3/U72/Z_26 , 
        \U3/U72/Z_25 , \U3/U72/Z_24 , \U3/U72/Z_23 , \U3/U72/Z_22 , 
        \U3/U72/Z_21 , \U3/U72/Z_20 , \U3/U72/Z_19 , \U3/U72/Z_18 , 
        \U3/U72/Z_17 , \U3/U72/Z_16 , \U3/U72/Z_15 , N2823, N2822, N2821, 
        N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, 
        N2810, N2417}), .B({\U3/U73/Z_31 , \U3/U73/Z_30 , \U3/U73/Z_29 , 
        \U3/U73/Z_28 , \U3/U73/Z_27 , \U3/U73/Z_26 , \U3/U73/Z_25 , 
        \U3/U73/Z_24 , \U3/U73/Z_23 , \U3/U73/Z_22 , \U3/U73/Z_21 , 
        \U3/U73/Z_20 , \U3/U73/Z_19 , \U3/U73/Z_18 , \U3/U73/Z_17 , 
        \U3/U73/Z_16 , \U3/U73/Z_15 , N2894, N2893, N2892, N2891, N2890, N2889, 
        N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2481}), .CI(
        1'b0), .SUM({N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, 
        N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, 
        N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, 
        N2388, N2387, N2386, N2385}) );
  CannyEdge_DW01_add_16 add_6_root_add_160_24 ( .A({N1642, N1641, N1640, N1639, 
        N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, 
        N1628}), .B({N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, 
        N1664, N1663, N1662, N1661, N1660, N1659, N1658}), .CI(1'b0), .SUM({
        N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, 
        N1872, N1871, N1870, N1869, N1868}) );
  CannyEdge_DW01_add_17 add_13_root_add_160_24 ( .A({N1927, N1926, N1925, 
        N1924, N1923, N1922, N1921, N1920, N1919, N1918, N3093, N3092, N3091, 
        N3090, N3089}), .B({N1957, N1956, N1955, N1954, N1953, N1952, N1951, 
        N1950, N1949, N3194, N3193, N3192, N3191, N3190, N3189}), .CI(1'b0), 
        .SUM({N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, 
        N1663, N1662, N1661, N1660, N1659, N1658}) );
  CannyEdge_DW01_add_18 add_14_root_add_160_24 ( .A({N1867, N1866, N1865, 
        N1864, N1863, N1862, N1861, N1860, N1859, N1858, N3343, N3342, N3341, 
        N3340, N3359}), .B({1'b0, N1896, N1895, N1894, N1893, N1892, N1891, 
        N1890, N1889, N976, N975, N974, N973, N972, N971}), .CI(1'b0), .SUM({
        N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, 
        N1632, N1631, N1630, N1629, N1628}) );
  CannyEdge_DW01_addsub_5 add_20_root_add_160_24 ( .A({1'b0, N1506, N1505, 
        N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, 
        N1494, N1493}), .B({1'b0, N1536, N1535, N1534, N1533, N1532, N1531, 
        N1530, N1529, N1528, N1527, N1526, N1525, N1524, 1'b0}), .CI(1'b0), 
        .ADD_SUB(1'b0), .SUM({N1462, N1461, N1460, N1459, N1458, N1457, N1456, 
        N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448}) );
  CannyEdge_DW01_addsub_7 r1802 ( .A({\U3/U78/Z_31 , \U3/U78/Z_30 , 
        \U3/U78/Z_29 , \U3/U78/Z_28 , \U3/U78/Z_27 , \U3/U78/Z_26 , 
        \U3/U78/Z_25 , \U3/U78/Z_24 , \U3/U78/Z_23 , \U3/U78/Z_22 , 
        \U3/U78/Z_21 , \U3/U78/Z_20 , \U3/U78/Z_19 , \U3/U78/Z_18 , 
        \U3/U78/Z_17 , \U3/U78/Z_16 , \U3/U78/Z_15 , \U3/U78/Z_14 , 
        \U3/U78/Z_13 , \U3/U78/Z_12 , \U3/U78/Z_11 , \U3/U78/Z_10 , 
        \U3/U78/Z_9 , \U3/U78/Z_8 , \U3/U78/Z_7 , \U3/U78/Z_6 , \U3/U78/Z_5 , 
        \U3/U78/Z_4 , \U3/U78/Z_3 , \U3/U78/Z_2 , \U3/U78/Z_1 , \U3/U78/Z_0 }), 
        .B({\U3/U79/Z_31 , \U3/U79/Z_30 , \U3/U79/Z_29 , \U3/U79/Z_28 , 
        \U3/U79/Z_27 , \U3/U79/Z_26 , \U3/U79/Z_25 , \U3/U79/Z_24 , 
        \U3/U79/Z_23 , \U3/U79/Z_22 , \U3/U79/Z_21 , \U3/U79/Z_20 , 
        \U3/U79/Z_19 , \U3/U79/Z_18 , \U3/U79/Z_17 , \U3/U79/Z_16 , 
        \U3/U79/Z_15 , \U3/U79/Z_14 , \U3/U79/Z_13 , \U3/U79/Z_12 , 
        \U3/U79/Z_11 , \U3/U79/Z_10 , \U3/U79/Z_9 , \U3/U79/Z_8 , \U3/U79/Z_7 , 
        \U3/U79/Z_6 , \U3/U79/Z_5 , \U3/U79/Z_4 , \U3/U79/Z_3 , \U3/U79/Z_2 , 
        \U3/U79/Z_1 , \U3/U79/Z_0 }), .CI(1'b0), .ADD_SUB(n7241), .SUM({N2331, 
        N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, 
        N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, 
        N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, 
        N2300}) );
  CannyEdge_DW01_add_19 add_1_root_add_202_8 ( .A({N2139, N2138, N2137, N2136, 
        N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, 
        N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, 
        N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108}), .B({N2203, 
        N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, 
        N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, 
        N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, 
        N2172}), .CI(1'b0), .SUM({N2299, N2298, N2297, N2296, N2295, N2294, 
        N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, 
        N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, 
        N2273, N2272, N2271, N2270, N2269, N2268}) );
  CannyEdge_DW01_add_20 r1223 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \U3/U70/Z_8 , \U3/U70/Z_7 , \U3/U70/Z_6 , 
        \U3/U70/Z_5 , \U3/U70/Z_4 , \U3/U70/Z_3 , \U3/U70/Z_2 , \U3/U70/Z_1 , 
        \U3/U70/Z_0 }), .B({\U3/U71/Z_31 , \U3/U71/Z_30 , \U3/U71/Z_29 , 
        \U3/U71/Z_28 , \U3/U71/Z_27 , \U3/U71/Z_26 , \U3/U71/Z_25 , 
        \U3/U71/Z_24 , \U3/U71/Z_23 , \U3/U71/Z_22 , \U3/U71/Z_21 , 
        \U3/U71/Z_20 , \U3/U71/Z_19 , \U3/U71/Z_18 , \U3/U71/Z_17 , 
        \U3/U71/Z_16 , \U3/U71/Z_15 , N2154, N2153, N2152, N2151, N2150, N2149, 
        N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140}), .CI(
        1'b0), .SUM({N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, 
        N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, 
        N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, 
        N2175, N2174, N2173, N2172}) );
  CannyEdge_DW01_add_21 r1814 ( .A({\U3/U68/Z_31 , \U3/U68/Z_30 , 
        \U3/U68/Z_29 , \U3/U68/Z_28 , \U3/U68/Z_27 , \U3/U68/Z_26 , 
        \U3/U68/Z_25 , \U3/U68/Z_24 , \U3/U68/Z_23 , \U3/U68/Z_22 , 
        \U3/U68/Z_21 , \U3/U68/Z_20 , \U3/U68/Z_19 , \U3/U68/Z_18 , 
        \U3/U68/Z_17 , \U3/U68/Z_16 , \U3/U68/Z_15 , N2090, N2089, N2088, 
        N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, 
        N2077, N2076}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U69/Z_13 , \U3/U69/Z_12 , \U3/U69/Z_11 , \U3/U69/Z_10 , 
        \U3/U69/Z_9 , \U3/U69/Z_8 , \U3/U69/Z_7 , \U3/U69/Z_6 , \U3/U69/Z_5 , 
        \U3/U69/Z_4 , \U3/U69/Z_3 , \U3/U69/Z_2 , \U3/U69/Z_1 , \U3/U69/Z_0 }), 
        .CI(1'b0), .SUM({N2139, N2138, N2137, N2136, N2135, N2134, N2133, 
        N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, 
        N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, 
        N2112, N2111, N2110, N2109, N2108}) );
  CannyEdge_DW01_addsub_9 r1201 ( .A({\U3/U100/Z_6 , n7203, n3691, n3692, 
        n3693, n3694, n3695}), .B({\U3/U101/Z_6 , \U3/U101/Z_6 , \U3/U101/Z_6 , 
        \U3/U101/Z_3 , n3690, n3689, \U3/U101/Z_0 }), .CI(1'b0), .ADD_SUB(1'b0), .SUM({N983, N982, N981, N980, N979, N978, N977}) );
  CannyEdge_DW01_addsub_11 r1337 ( .A({\U3/U134/Z_10 , \U3/U134/Z_9 , 
        \U3/U134/Z_8 , \U3/U134/Z_7 , \U3/U134/Z_6 , \U3/U134/Z_5 , 
        \U3/U134/Z_4 , \U3/U134/Z_3 , \U3/U134/Z_2 , \U3/U134/Z_1 , 
        \U3/U134/Z_0 }), .B({n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
        n3703, n3704, n3705, n3706}), .CI(1'b0), .ADD_SUB(\U3/U136/Z_0 ), 
        .SUM({N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  CannyEdge_DW01_addsub_12 r1343 ( .A(Gx[10:0]), .B(Gy[10:0]), .CI(1'b0), 
        .ADD_SUB(n3707), .SUM({N2568, N2567, N2566, N2565, N2564, N2563, N2562, 
        N2561, N2560, N2559, N2558}) );
  CannyEdge_DW01_cmp2_0 lte_289 ( .A(fGy), .B({N2840, N2840, N2839, N2838, 
        N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, 
        N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, 
        N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810}), .LEQ(1'b1), 
        .TC(1'b1), .LT_LE(N2841) );
  CannyEdge_DW01_cmp2_1 gt_274 ( .A({N2911, N2911, N2910, N2909, N2908, N2907, 
        N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, 
        N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, 
        N2886, N2885, N2884, N2883, N2882, N2881}), .B(fGy), .LEQ(1'b0), .TC(
        1'b1), .LT_LE(N2945) );
  CannyEdge_DW01_cmp2_2 gt_292 ( .A({N2840, N2840, N2839, N2838, N2837, N2836, 
        N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, 
        N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, 
        N2815, N2814, N2813, N2812, N2811, N2810}), .B(fGy), .LEQ(1'b0), .TC(
        1'b1), .LT_LE(N2874) );
  CannyEdge_DW02_mult_0 mult_160_18 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[17][7] , \regX[17][6] , \regX[17][5] , 
        \regX[17][4] , \regX[17][3] , \regX[17][2] , \regX[17][1] , 
        \regX[17][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, N1836, N1835, N1834, N1833, N1832, N1831, 
        N1830, N1829, N1828, N1827, N1826, N1825, N1824, 
        SYNOPSYS_UNCONNECTED__13}) );
  CannyEdge_DW02_mult_1 mult_160_17 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[16][7] , \regX[16][6] , \regX[16][5] , 
        \regX[16][4] , \regX[16][3] , \regX[16][2] , \regX[16][1] , 
        \regX[16][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N1806, N1805, N1804, N1803, N1802, N1801, 
        N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793}) );
  CannyEdge_DW02_mult_2 mult_160_16 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[15][7] , \regX[15][6] , \regX[15][5] , 
        \regX[15][4] , \regX[15][3] , \regX[15][2] , \regX[15][1] , 
        \regX[15][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, N1776, N1775, N1774, N1773, N1772, N1771, 
        N1770, N1769, N1768, N1767, N1766, N1765, N1569, N1568}) );
  CannyEdge_DW02_mult_4 mult_160_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[13][7] , \regX[13][6] , \regX[13][5] , 
        \regX[13][4] , \regX[13][3] , \regX[13][2] , \regX[13][1] , 
        \regX[13][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, N1716, N1715, N1714, N1713, N1712, N1711, 
        N1710, N1709, N1708, N1707, N1541, N1540, N1539, 
        SYNOPSYS_UNCONNECTED__20}) );
  CannyEdge_DW02_mult_6 mult_160_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[11][7] , \regX[11][6] , \regX[11][5] , 
        \regX[11][4] , \regX[11][3] , \regX[11][2] , \regX[11][1] , 
        \regX[11][0] }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, N1656, N1655, N1654, N1653, N1652, N1651, 
        N1650, N1649, N1648, N1647, N1646, N1645, N1509, 
        SYNOPSYS_UNCONNECTED__23}) );
  CannyEdge_DW02_mult_8 mult_160_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[9][7] , \regX[9][6] , \regX[9][5] , 
        \regX[9][4] , \regX[9][3] , \regX[9][2] , \regX[9][1] , \regX[9][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, N1596, N1595, N1594, N1593, N1592, N1591, 
        N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583}) );
  CannyEdge_DW02_mult_9 mult_160_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[8][7] , \regX[8][6] , \regX[8][5] , 
        \regX[8][4] , \regX[8][3] , \regX[8][2] , \regX[8][1] , \regX[8][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N1566, N1565, N1564, N1563, N1562, N1561, 
        N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553}) );
  CannyEdge_DW02_mult_10 mult_160_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0}), .B({\regX[7][7] , \regX[7][6] , \regX[7][5] , 
        \regX[7][4] , \regX[7][3] , \regX[7][2] , \regX[7][1] , \regX[7][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, N1536, N1535, N1534, N1533, N1532, N1531, 
        N1530, N1529, N1528, N1527, N1526, N1525, N1524, 
        SYNOPSYS_UNCONNECTED__30}) );
  CannyEdge_DW02_mult_11 r1229 ( .A({n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n3484, n3483, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n2980, n7253}), .B({\regX[5][7] , 
        \regX[5][6] , \regX[5][5] , \regX[5][4] , \regX[5][3] , \regX[5][2] , 
        \regX[5][1] , \regX[5][0] }), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, N2171, N2170, 
        N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, 
        N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, 
        N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140})
         );
  CannyEdge_DW02_mult_14 mult_160_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b1}), .B({\regX[1][7] , \regX[1][6] , \regX[1][5] , 
        \regX[1][4] , \regX[1][3] , \regX[1][2] , \regX[1][1] , \regX[1][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, N1356, N1355, N1354, N1353, N1352, N1351, 
        N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343}) );
  CannyEdge_DW02_mult_15 r1211 ( .A({n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n3484, n3483, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n2980}), .B({\regX[0][7] , 
        \regX[0][6] , \regX[0][5] , \regX[0][4] , \regX[0][3] , \regX[0][2] , 
        \regX[0][1] , \regX[0][0] }), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, N2107, N2106, 
        N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, 
        N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, 
        N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076})
         );
  CannyEdge_DW02_mult_16 r1207 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n4572, 
        n4573, n4574}), .B({\U3/U63/Z_7 , \U3/U63/Z_6 , \U3/U63/Z_5 , 
        \U3/U63/Z_4 , \U3/U63/Z_3 , \U3/U63/Z_2 , \U3/U63/Z_1 , \U3/U63/Z_0 }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, N1896, N1895, N1894, N1893, N1892, N1891, 
        N1890, N1889, N976, N975, N974, N973, N972, N971}) );
  CannyEdge_DW02_mult_17 r1075 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n7202, 
        n7253, \U3/U124/Z_0 }), .B({\U3/U125/Z_7 , \U3/U125/Z_6 , 
        \U3/U125/Z_5 , \U3/U125/Z_4 , \U3/U125/Z_3 , \U3/U125/Z_2 , 
        \U3/U125/Z_1 , \U3/U125/Z_0 }), .TC(n7202), .PRODUCT({
        SYNOPSYS_UNCONNECTED__51, N1417, N1416, N1415, N1414, N1413, N1412, 
        N1411, N1410, N1409, N1408, N3443, N3442, N3441, N1389, N1388}) );
  CannyEdge_DW02_mult_18 r1062 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n7204, 
        n7253, \U3/U97/Z_0 }), .B({\U3/U98/Z_7 , \U3/U98/Z_6 , \U3/U98/Z_5 , 
        \U3/U98/Z_4 , \U3/U98/Z_3 , \U3/U98/Z_2 , \U3/U98/Z_1 , \U3/U98/Z_0 }), 
        .TC(n7204), .PRODUCT({SYNOPSYS_UNCONNECTED__52, N1957, N1956, N1955, 
        N1954, N1953, N1952, N1951, N1950, N1949, N3194, N3193, N3192, N3191, 
        N3190, N3189}) );
  CannyEdge_DW01_cmp2_3 r1050 ( .A({n7211, n7212, n7213, n7214, n7215, n7216, 
        n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, 
        n7227, n7228, n7229, n7230, n7231, n7232, n7209, n7210, \U3/U121/Z_7 , 
        \U3/U121/Z_6 , \U3/U121/Z_5 , \U3/U121/Z_4 , \U3/U121/Z_3 , 
        \U3/U121/Z_2 , \U3/U121/Z_1 , \U3/U121/Z_0 }), .B({1'b0, 1'b0, 
        \U3/U122/Z_29 , \U3/U122/Z_28 , \U3/U122/Z_27 , \U3/U122/Z_26 , 
        \U3/U122/Z_25 , \U3/U122/Z_24 , \U3/U122/Z_23 , \U3/U122/Z_22 , 
        \U3/U122/Z_21 , \U3/U122/Z_20 , \U3/U122/Z_19 , \U3/U122/Z_18 , 
        \U3/U122/Z_17 , \U3/U122/Z_16 , \U3/U122/Z_15 , \U3/U122/Z_14 , 
        \U3/U122/Z_13 , \U3/U122/Z_12 , \U3/U122/Z_11 , \U3/U122/Z_10 , 
        \U3/U122/Z_9 , \U3/U122/Z_8 , \U3/U122/Z_7 , \U3/U122/Z_6 , 
        \U3/U122/Z_5 , \U3/U122/Z_4 , \U3/U122/Z_3 , \U3/U122/Z_2 , 
        \U3/U122/Z_1 , \U3/U122/Z_0 }), .LEQ(1'b1), .TC(n7240), .GE_GT(N2880)
         );
  CannyEdge_DW02_mult_19 r1047 ( .A({\U3/U84/Z_7 , \U3/U84/Z_6 , \U3/U84/Z_5 , 
        \U3/U84/Z_4 , \U3/U84/Z_3 , \U3/U84/Z_2 , \U3/U84/Z_1 , \U3/U84/Z_0 }), 
        .B({\U3/U85/Z_31 , \U3/U85/Z_30 , \U3/U85/Z_29 , \U3/U85/Z_28 , 
        \U3/U85/Z_27 , \U3/U85/Z_26 , \U3/U85/Z_25 , \U3/U85/Z_24 , 
        \U3/U85/Z_23 , \U3/U85/Z_22 , \U3/U85/Z_21 , \U3/U85/Z_20 , 
        \U3/U85/Z_19 , \U3/U85/Z_18 , \U3/U85/Z_17 , \U3/U85/Z_16 , 
        \U3/U85/Z_15 , \U3/U85/Z_14 , \U3/U85/Z_13 , \U3/U85/Z_12 , 
        \U3/U85/Z_11 , \U3/U85/Z_10 , \U3/U85/Z_9 , \U3/U85/Z_8 , \U3/U85/Z_7 , 
        \U3/U85/Z_6 , \U3/U85/Z_5 , \U3/U85/Z_4 , \U3/U85/Z_3 , \U3/U85/Z_2 , 
        \U3/U85/Z_1 , \U3/U85/Z_0 }), .TC(n3467), .PRODUCT({
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, N2840, N2839, 
        N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, 
        N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, 
        N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2417})
         );
  CannyEdge_DW01_cmp2_4 r1033 ( .A({\U3/U93/Z_31 , \U3/U93/Z_30 , 
        \U3/U93/Z_29 , \U3/U93/Z_28 , \U3/U93/Z_27 , \U3/U93/Z_26 , 
        \U3/U93/Z_25 , \U3/U93/Z_24 , \U3/U93/Z_23 , \U3/U93/Z_22 , 
        \U3/U93/Z_21 , \U3/U93/Z_20 , \U3/U93/Z_19 , \U3/U93/Z_18 , 
        \U3/U93/Z_17 , \U3/U93/Z_16 , \U3/U93/Z_15 , \U3/U93/Z_14 , 
        \U3/U93/Z_13 , \U3/U93/Z_12 , \U3/U93/Z_11 , \U3/U93/Z_10 , 
        \U3/U93/Z_9 , \U3/U93/Z_8 , \U3/U93/Z_7 , \U3/U93/Z_6 , \U3/U93/Z_5 , 
        \U3/U93/Z_4 , \U3/U93/Z_3 , \U3/U93/Z_2 , \U3/U93/Z_1 , \U3/U93/Z_0 }), 
        .B({\U3/U94/Z_31 , \U3/U94/Z_31 , \U3/U94/Z_29 , \U3/U94/Z_28 , 
        \U3/U94/Z_27 , \U3/U94/Z_26 , \U3/U94/Z_25 , \U3/U94/Z_24 , 
        \U3/U94/Z_23 , \U3/U94/Z_22 , \U3/U94/Z_21 , \U3/U94/Z_20 , 
        \U3/U94/Z_19 , \U3/U94/Z_18 , \U3/U94/Z_17 , \U3/U94/Z_16 , 
        \U3/U94/Z_15 , \U3/U94/Z_14 , \U3/U94/Z_13 , \U3/U94/Z_12 , 
        \U3/U94/Z_11 , \U3/U94/Z_10 , \U3/U94/Z_9 , \U3/U94/Z_8 , \U3/U94/Z_7 , 
        \U3/U94/Z_6 , \U3/U94/Z_5 , \U3/U94/Z_4 , \U3/U94/Z_3 , \U3/U94/Z_2 , 
        \U3/U94/Z_1 , \U3/U94/Z_0 }), .LEQ(\U3/U95/Z_0 ), .TC(\U3/U96/Z_0 ), 
        .GE_GT(N2549) );
  CannyEdge_DW02_mult_20 r1051 ( .A({\U3/U87/Z_7 , \U3/U87/Z_6 , \U3/U87/Z_5 , 
        \U3/U87/Z_4 , \U3/U87/Z_3 , \U3/U87/Z_2 , \U3/U87/Z_1 , \U3/U87/Z_0 }), 
        .B({n3483, \U3/U88/Z_30 , \U3/U88/Z_29 , \U3/U88/Z_28 , \U3/U88/Z_27 , 
        \U3/U88/Z_26 , \U3/U88/Z_25 , \U3/U88/Z_24 , \U3/U88/Z_23 , 
        \U3/U88/Z_22 , \U3/U88/Z_21 , \U3/U88/Z_20 , \U3/U88/Z_19 , 
        \U3/U88/Z_18 , \U3/U88/Z_17 , \U3/U88/Z_16 , \U3/U88/Z_15 , 
        \U3/U88/Z_14 , \U3/U88/Z_13 , \U3/U88/Z_12 , \U3/U88/Z_11 , 
        \U3/U88/Z_10 , \U3/U88/Z_9 , \U3/U88/Z_8 , \U3/U88/Z_7 , \U3/U88/Z_6 , 
        \U3/U88/Z_5 , \U3/U88/Z_4 , \U3/U88/Z_3 , \U3/U88/Z_2 , \U3/U88/Z_1 , 
        \U3/U88/Z_0 }), .TC(n7240), .PRODUCT({SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, N2911, N2910, N2909, N2908, N2907, N2906, 
        N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, 
        N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, 
        N2885, N2884, N2883, N2882, N2881, N2481}) );
  CannyEdge_DW02_mult_21 mult_160_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b1, 1'b1}), .B({\regX[6][7] , \regX[6][6] , \regX[6][5] , 
        \regX[6][4] , \regX[6][3] , \regX[6][2] , \regX[6][1] , \regX[6][0] }), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, N1506, N1505, N1504, N1503, N1502, N1501, 
        N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493}) );
  CannyEdge_DW01_cmp2_5 r169 ( .A({\U3/U118/Z_31 , \U3/U118/Z_30 , 
        \U3/U118/Z_29 , \U3/U118/Z_28 , \U3/U118/Z_27 , \U3/U118/Z_26 , 
        \U3/U118/Z_25 , \U3/U118/Z_24 , \U3/U118/Z_23 , \U3/U118/Z_22 , 
        \U3/U118/Z_21 , \U3/U118/Z_20 , \U3/U118/Z_19 , \U3/U118/Z_18 , 
        \U3/U118/Z_17 , \U3/U118/Z_16 , \U3/U118/Z_15 , \U3/U118/Z_14 , 
        \U3/U118/Z_13 , \U3/U118/Z_12 , \U3/U118/Z_11 , \U3/U118/Z_10 , 
        \U3/U118/Z_9 , \U3/U118/Z_8 , \U3/U118/Z_7 , \U3/U118/Z_6 , 
        \U3/U118/Z_5 , \U3/U118/Z_4 , \U3/U118/Z_3 , \U3/U118/Z_2 , 
        \U3/U118/Z_1 , \U3/U118/Z_0 }), .B({\U3/U119/Z_31 , \U3/U119/Z_31 , 
        \U3/U119/Z_29 , \U3/U119/Z_28 , \U3/U119/Z_27 , \U3/U119/Z_26 , 
        \U3/U119/Z_25 , \U3/U119/Z_24 , \U3/U119/Z_23 , \U3/U119/Z_22 , 
        \U3/U119/Z_21 , \U3/U119/Z_20 , \U3/U119/Z_19 , \U3/U119/Z_18 , 
        \U3/U119/Z_17 , \U3/U119/Z_16 , \U3/U119/Z_15 , \U3/U119/Z_14 , 
        \U3/U119/Z_13 , \U3/U119/Z_12 , \U3/U119/Z_11 , \U3/U119/Z_10 , 
        \U3/U119/Z_9 , \U3/U119/Z_8 , \U3/U119/Z_7 , \U3/U119/Z_6 , 
        \U3/U119/Z_5 , \U3/U119/Z_4 , \U3/U119/Z_3 , \U3/U119/Z_2 , 
        \U3/U119/Z_1 , \U3/U119/Z_0 }), .LEQ(1'b1), .TC(n3467), .LT_LE(N2777)
         );
  CannyEdge_DW02_mult_22 r1055 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n7246, 1'b0, 
        \U3/U90/Z_0 }), .B({\U3/U91/Z_7 , \U3/U91/Z_6 , \U3/U91/Z_5 , 
        \U3/U91/Z_4 , \U3/U91/Z_3 , \U3/U91/Z_2 , \U3/U91/Z_1 , \U3/U91/Z_0 }), 
        .TC(n7246), .PRODUCT({SYNOPSYS_UNCONNECTED__71, N1927, N1926, N1925, 
        N1924, N1923, N1922, N1921, N1920, N1919, N1918, N3093, N3092, N3091, 
        N3090, N3089}) );
  CannyEdge_DW02_mult_23 r1068 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \U3/U109/Z_2 , n7253, \U3/U109/Z_2 }), .B({\U3/U110/Z_7 , 
        \U3/U110/Z_6 , \U3/U110/Z_5 , \U3/U110/Z_4 , \U3/U110/Z_3 , 
        \U3/U110/Z_2 , \U3/U110/Z_1 , \U3/U110/Z_0 }), .TC(n7205), .PRODUCT({
        SYNOPSYS_UNCONNECTED__72, N1867, N1866, N1865, N1864, N1863, N1862, 
        N1861, N1860, N1859, N1858, N3343, N3342, N3341, N3340, N3359}) );
  CannyEdge_DW01_cmp2_6 r1377 ( .A({\U3/U119/Z_31 , \U3/U119/Z_31 , 
        \U3/U119/Z_29 , \U3/U119/Z_28 , \U3/U119/Z_27 , \U3/U119/Z_26 , 
        \U3/U119/Z_25 , \U3/U119/Z_24 , \U3/U119/Z_23 , \U3/U119/Z_22 , 
        \U3/U119/Z_21 , \U3/U119/Z_20 , \U3/U119/Z_19 , \U3/U119/Z_18 , 
        \U3/U119/Z_17 , \U3/U119/Z_16 , \U3/U119/Z_15 , \U3/U119/Z_14 , 
        \U3/U119/Z_13 , \U3/U119/Z_12 , \U3/U119/Z_11 , \U3/U119/Z_10 , 
        \U3/U119/Z_9 , \U3/U119/Z_8 , n7242, n7243, n7244, n7245, 
        \U3/U105/Z_3 , \U3/U105/Z_2 , \U3/U105/Z_1 , \U3/U105/Z_0 }), .B({
        \U3/U118/Z_31 , \U3/U118/Z_30 , \U3/U118/Z_29 , \U3/U118/Z_28 , 
        \U3/U118/Z_27 , \U3/U118/Z_26 , \U3/U118/Z_25 , \U3/U118/Z_24 , 
        \U3/U118/Z_23 , \U3/U118/Z_22 , \U3/U118/Z_21 , \U3/U118/Z_20 , 
        \U3/U118/Z_19 , \U3/U118/Z_18 , \U3/U118/Z_17 , \U3/U118/Z_16 , 
        \U3/U118/Z_15 , \U3/U118/Z_14 , \U3/U118/Z_13 , \U3/U118/Z_12 , 
        \U3/U118/Z_11 , \U3/U118/Z_10 , \U3/U118/Z_9 , \U3/U118/Z_8 , n7247, 
        n7248, n7249, n7250, \U3/U106/Z_3 , n7251, \U3/U106/Z_1 , n7252}), 
        .LEQ(n4612), .TC(n3467), .LT_LE(N3336) );
  CannyEdge_DW01_addsub_16 r1044 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \U3/U81/Z_7 , \U3/U81/Z_6 , 
        \U3/U81/Z_5 , \U3/U81/Z_4 , \U3/U81/Z_3 , \U3/U81/Z_2 , \U3/U81/Z_1 , 
        \U3/U81/Z_0 }), .B({\U3/U82/Z_31 , \U3/U82/Z_30 , \U3/U82/Z_29 , 
        \U3/U82/Z_28 , \U3/U82/Z_27 , \U3/U82/Z_26 , \U3/U82/Z_25 , 
        \U3/U82/Z_24 , \U3/U82/Z_23 , \U3/U82/Z_22 , \U3/U82/Z_21 , 
        \U3/U82/Z_20 , \U3/U82/Z_19 , \U3/U82/Z_18 , \U3/U82/Z_17 , 
        \U3/U82/Z_16 , \U3/U82/Z_15 , \U3/U82/Z_14 , \U3/U82/Z_13 , 
        \U3/U82/Z_12 , \U3/U82/Z_11 , \U3/U82/Z_10 , \U3/U82/Z_9 , 
        \U3/U82/Z_8 , \U3/U82/Z_7 , \U3/U82/Z_6 , \U3/U82/Z_5 , \U3/U82/Z_4 , 
        \U3/U82/Z_3 , \U3/U82/Z_2 , \U3/U82/Z_1 , \U3/U82/Z_0 }), .CI(1'b0), 
        .ADD_SUB(n3473), .SUM({N2776, N2775, N2774, N2773, N2772, N2771, N2770, 
        N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, 
        N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, 
        N2749, N2748, N2747, N2746, N2648}) );
  CannyEdge_DW02_mult_24 r1023 ( .A({\U3/U64/Z_7 , \U3/U64/Z_6 , \U3/U64/Z_5 , 
        \U3/U64/Z_4 , \U3/U64/Z_3 , \U3/U64/Z_2 , \U3/U64/Z_1 , \U3/U64/Z_0 }), 
        .B({n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, n3484, 
        n3484, n3484, n3484, n3483, n3484, \U3/U65/Z_7 , \U3/U65/Z_6 , 
        \U3/U65/Z_5 , \U3/U65/Z_4 , \U3/U65/Z_3 , \U3/U65/Z_2 , \U3/U65/Z_1 , 
        \U3/U65/Z_0 }), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, N2267, N2266, N2265, N2264, N2263, N2262, 
        N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, 
        N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, 
        N2241, N2240, N2239, N2238, N2237, N2236}) );
  AND2X2 U23 ( .A(n5457), .B(n4131), .Y(n3467) );
  OR2X2 U26 ( .A(n3488), .B(n3471), .Y(n3468) );
  AND2X2 U27 ( .A(n4127), .B(n4128), .Y(n3469) );
  AND2X2 U28 ( .A(n3480), .B(n3471), .Y(n3470) );
  INVX2 U29 ( .A(n3469), .Y(n3471) );
  INVX2 U30 ( .A(n3468), .Y(n3472) );
  INVX4 U32 ( .A(n3470), .Y(n3473) );
  INVX4 U35 ( .A(n5790), .Y(n3946) );
  INVX1 U36 ( .A(n5823), .Y(n3474) );
  INVX4 U37 ( .A(n3474), .Y(n3475) );
  INVX4 U38 ( .A(n3488), .Y(n3555) );
  INVX4 U39 ( .A(n3484), .Y(n3476) );
  INVX4 U40 ( .A(n3467), .Y(n3477) );
  INVX2 U41 ( .A(n3949), .Y(n3478) );
  INVX2 U42 ( .A(n5827), .Y(n7246) );
  INVX2 U43 ( .A(n4257), .Y(n3479) );
  INVX4 U44 ( .A(n3548), .Y(n4257) );
  INVX2 U45 ( .A(n5457), .Y(n3480) );
  BUFX2 U46 ( .A(n3552), .Y(n3481) );
  AND2X2 U47 ( .A(n4015), .B(n4127), .Y(n4025) );
  INVX2 U49 ( .A(n7240), .Y(n3482) );
  INVX2 U51 ( .A(n5826), .Y(n7240) );
  INVX2 U52 ( .A(n3475), .Y(n7253) );
  INVX4 U53 ( .A(n3471), .Y(n7241) );
  INVX4 U56 ( .A(n5791), .Y(n3483) );
  INVX2 U59 ( .A(n5791), .Y(n3484) );
  INVX1 U61 ( .A(n3485), .Y(n7200) );
  MUX2X1 U63 ( .B(\regY[6][6] ), .A(InData[6]), .S(n3486), .Y(n3485) );
  INVX1 U64 ( .A(n3487), .Y(n7201) );
  AOI22X1 U65 ( .A(n3488), .B(fGy[31]), .C(n3472), .D(N2776), .Y(n3487) );
  INVX1 U66 ( .A(n3489), .Y(n7203) );
  AOI21X1 U67 ( .A(n3490), .B(N976), .C(\U3/U100/Z_6 ), .Y(n3489) );
  INVX1 U68 ( .A(n3491), .Y(n7206) );
  AOI22X1 U69 ( .A(N2341), .B(n3483), .C(N2394), .D(n7253), .Y(n3491) );
  INVX1 U70 ( .A(n3492), .Y(n7207) );
  AOI22X1 U72 ( .A(N2340), .B(n3483), .C(N2393), .D(n7253), .Y(n3492) );
  INVX1 U74 ( .A(n3493), .Y(n7208) );
  AOI22X1 U76 ( .A(N2339), .B(n3483), .C(N2392), .D(n7253), .Y(n3493) );
  INVX1 U77 ( .A(n3494), .Y(n7209) );
  INVX1 U78 ( .A(n3495), .Y(n7210) );
  INVX1 U79 ( .A(n3496), .Y(n7211) );
  INVX1 U82 ( .A(n3497), .Y(n7212) );
  INVX1 U83 ( .A(n3498), .Y(n7213) );
  INVX1 U84 ( .A(n3499), .Y(n7214) );
  INVX1 U90 ( .A(n3500), .Y(n7215) );
  INVX1 U97 ( .A(n3501), .Y(n7216) );
  INVX1 U99 ( .A(n3502), .Y(n7217) );
  INVX1 U114 ( .A(n3503), .Y(n7218) );
  INVX1 U116 ( .A(n3504), .Y(n7219) );
  INVX1 U210 ( .A(n3505), .Y(n7220) );
  INVX1 U211 ( .A(n3506), .Y(n7221) );
  INVX1 U212 ( .A(n3507), .Y(n7222) );
  INVX1 U213 ( .A(n3508), .Y(n7223) );
  INVX1 U214 ( .A(n3509), .Y(n7224) );
  INVX1 U215 ( .A(n3510), .Y(n7225) );
  INVX1 U216 ( .A(n3511), .Y(n7226) );
  INVX1 U217 ( .A(n3512), .Y(n7227) );
  INVX1 U218 ( .A(n3513), .Y(n7228) );
  INVX1 U219 ( .A(n3514), .Y(n7229) );
  INVX1 U220 ( .A(n3515), .Y(n7230) );
  INVX1 U221 ( .A(n3516), .Y(n7231) );
  INVX1 U222 ( .A(n3517), .Y(n7232) );
  INVX1 U223 ( .A(n3518), .Y(n7233) );
  AOI22X1 U224 ( .A(N2338), .B(n3483), .C(N2391), .D(n7253), .Y(n3518) );
  INVX1 U225 ( .A(n3519), .Y(n7234) );
  AOI22X1 U226 ( .A(N2337), .B(n3483), .C(N2390), .D(n7253), .Y(n3519) );
  INVX1 U227 ( .A(n3520), .Y(n7235) );
  AOI22X1 U228 ( .A(N2336), .B(n3483), .C(N2389), .D(n7253), .Y(n3520) );
  INVX1 U229 ( .A(n3521), .Y(n7236) );
  AOI22X1 U230 ( .A(N2335), .B(n3483), .C(N2388), .D(n7253), .Y(n3521) );
  INVX1 U231 ( .A(n3522), .Y(n7237) );
  AOI22X1 U232 ( .A(N2334), .B(n3483), .C(N2387), .D(n7253), .Y(n3522) );
  INVX1 U233 ( .A(n3523), .Y(n7238) );
  AOI22X1 U234 ( .A(N2333), .B(n3483), .C(N2386), .D(n7253), .Y(n3523) );
  INVX1 U235 ( .A(n3524), .Y(n7239) );
  AOI22X1 U236 ( .A(N2332), .B(n3483), .C(N2385), .D(n7253), .Y(n3524) );
  INVX1 U237 ( .A(n3525), .Y(n7242) );
  INVX1 U238 ( .A(n3526), .Y(n7243) );
  INVX1 U239 ( .A(n3527), .Y(n7244) );
  INVX1 U240 ( .A(n3528), .Y(n7245) );
  INVX1 U241 ( .A(n3529), .Y(n7247) );
  INVX1 U242 ( .A(n3530), .Y(n7248) );
  INVX1 U243 ( .A(n3531), .Y(n7249) );
  INVX1 U244 ( .A(n3532), .Y(n7250) );
  INVX1 U245 ( .A(n3533), .Y(n7251) );
  INVX1 U246 ( .A(n3534), .Y(n7252) );
  INVX1 U247 ( .A(N4468), .Y(n7730) );
  INVX1 U248 ( .A(N4471), .Y(n7731) );
  INVX1 U249 ( .A(N4474), .Y(n7732) );
  INVX1 U250 ( .A(N4477), .Y(n7733) );
  INVX1 U251 ( .A(N4480), .Y(n7734) );
  INVX1 U252 ( .A(N4483), .Y(n7735) );
  INVX1 U253 ( .A(N4486), .Y(n7736) );
  OAI21X1 U254 ( .A(n7254), .B(n3535), .C(n3536), .Y(n5443) );
  INVX1 U255 ( .A(N4469), .Y(n7254) );
  OAI21X1 U256 ( .A(n7255), .B(n3535), .C(n3536), .Y(n5442) );
  INVX1 U257 ( .A(N4472), .Y(n7255) );
  OAI21X1 U258 ( .A(n7256), .B(n3535), .C(n3536), .Y(n5441) );
  INVX1 U259 ( .A(N4475), .Y(n7256) );
  OAI21X1 U260 ( .A(n7257), .B(n3535), .C(n3536), .Y(n5440) );
  INVX1 U261 ( .A(N4478), .Y(n7257) );
  OAI21X1 U262 ( .A(n7258), .B(n3535), .C(n3536), .Y(n5439) );
  INVX1 U263 ( .A(N4481), .Y(n7258) );
  OAI21X1 U264 ( .A(n7259), .B(n3535), .C(n3536), .Y(n5438) );
  INVX1 U265 ( .A(N4484), .Y(n7259) );
  OAI21X1 U266 ( .A(n7260), .B(n3535), .C(n3536), .Y(n5437) );
  INVX1 U267 ( .A(N4487), .Y(n7260) );
  OAI21X1 U268 ( .A(n7261), .B(n3535), .C(n3536), .Y(n5436) );
  NAND3X1 U269 ( .A(n3537), .B(n3538), .C(n3535), .Y(n3536) );
  INVX1 U270 ( .A(n3539), .Y(n3538) );
  INVX1 U271 ( .A(N4490), .Y(n7261) );
  OAI21X1 U272 ( .A(n3540), .B(n3541), .C(n3542), .Y(n5435) );
  OAI21X1 U273 ( .A(n3543), .B(n3544), .C(n3545), .Y(n3542) );
  OAI22X1 U274 ( .A(n3546), .B(n3547), .C(n3548), .D(n3549), .Y(n3544) );
  OR2X1 U275 ( .A(n3467), .B(n2980), .Y(n3543) );
  OAI21X1 U276 ( .A(n3546), .B(n3550), .C(n3551), .Y(n3541) );
  OAI22X1 U277 ( .A(n3550), .B(n3481), .C(n3553), .D(n3554), .Y(n5434) );
  INVX1 U278 ( .A(n3551), .Y(n3553) );
  NAND2X1 U279 ( .A(bOPEnable), .B(bCE), .Y(n3551) );
  OAI21X1 U280 ( .A(n7262), .B(n3555), .C(n3556), .Y(n5433) );
  INVX1 U281 ( .A(N4394), .Y(n7262) );
  OAI21X1 U282 ( .A(n7263), .B(n3555), .C(n3556), .Y(n5432) );
  INVX1 U283 ( .A(N4391), .Y(n7263) );
  OAI21X1 U284 ( .A(n7264), .B(n3555), .C(n3556), .Y(n5431) );
  INVX1 U285 ( .A(N4388), .Y(n7264) );
  OAI21X1 U286 ( .A(n7265), .B(n3555), .C(n3556), .Y(n5430) );
  INVX1 U287 ( .A(N4385), .Y(n7265) );
  OAI21X1 U288 ( .A(n7266), .B(n3555), .C(n3556), .Y(n5429) );
  INVX1 U289 ( .A(N4382), .Y(n7266) );
  OAI21X1 U290 ( .A(n7267), .B(n3555), .C(n3556), .Y(n5428) );
  INVX1 U291 ( .A(N4379), .Y(n7267) );
  OAI21X1 U292 ( .A(n7268), .B(n3555), .C(n3556), .Y(n5427) );
  INVX1 U293 ( .A(N4376), .Y(n7268) );
  OAI21X1 U294 ( .A(n7269), .B(n3555), .C(n3556), .Y(n5426) );
  INVX1 U295 ( .A(N4373), .Y(n7269) );
  OAI21X1 U296 ( .A(n7270), .B(n3555), .C(n3556), .Y(n5425) );
  INVX1 U297 ( .A(N4466), .Y(n7270) );
  OAI21X1 U298 ( .A(n7271), .B(n3555), .C(n3556), .Y(n5424) );
  INVX1 U299 ( .A(N4463), .Y(n7271) );
  OAI21X1 U300 ( .A(n7272), .B(n3555), .C(n3556), .Y(n5423) );
  INVX1 U301 ( .A(N4460), .Y(n7272) );
  OAI21X1 U302 ( .A(n7273), .B(n3555), .C(n3556), .Y(n5422) );
  INVX1 U303 ( .A(N4457), .Y(n7273) );
  OAI21X1 U304 ( .A(n7274), .B(n3555), .C(n3556), .Y(n5421) );
  INVX1 U305 ( .A(N4454), .Y(n7274) );
  OAI21X1 U306 ( .A(n7275), .B(n3555), .C(n3556), .Y(n5420) );
  INVX1 U307 ( .A(N4451), .Y(n7275) );
  OAI21X1 U308 ( .A(n7276), .B(n3555), .C(n3556), .Y(n5419) );
  INVX1 U309 ( .A(N4448), .Y(n7276) );
  OAI21X1 U310 ( .A(n7277), .B(n3555), .C(n3556), .Y(n5418) );
  NAND2X1 U311 ( .A(n3557), .B(n3555), .Y(n3556) );
  INVX1 U312 ( .A(N4445), .Y(n7277) );
  OAI21X1 U313 ( .A(n7278), .B(n3558), .C(n3559), .Y(n5417) );
  INVX1 U314 ( .A(N4502), .Y(n7278) );
  MUX2X1 U315 ( .B(n3560), .A(n3561), .S(n3562), .Y(n5416) );
  MUX2X1 U316 ( .B(n3563), .A(n3564), .S(n3562), .Y(n5415) );
  MUX2X1 U317 ( .B(n3565), .A(n3566), .S(n3562), .Y(n5414) );
  MUX2X1 U318 ( .B(n3567), .A(n3568), .S(n3562), .Y(n5413) );
  MUX2X1 U319 ( .B(n3569), .A(n3570), .S(n3562), .Y(n5412) );
  MUX2X1 U320 ( .B(n3571), .A(n3572), .S(n3562), .Y(n5411) );
  MUX2X1 U321 ( .B(n3573), .A(n3574), .S(n3562), .Y(n5410) );
  MUX2X1 U322 ( .B(n3575), .A(n3576), .S(n3562), .Y(n5409) );
  OAI21X1 U323 ( .A(n3577), .B(n3578), .C(n3579), .Y(n3562) );
  NAND3X1 U324 ( .A(n3580), .B(n3581), .C(n3582), .Y(n3579) );
  NAND2X1 U325 ( .A(n3583), .B(n3584), .Y(n3578) );
  NAND2X1 U326 ( .A(n3585), .B(n3586), .Y(n3577) );
  MUX2X1 U327 ( .B(n3587), .A(n3561), .S(n3588), .Y(n5408) );
  MUX2X1 U328 ( .B(n3589), .A(n3564), .S(n3588), .Y(n5407) );
  MUX2X1 U329 ( .B(n3590), .A(n3566), .S(n3588), .Y(n5406) );
  MUX2X1 U330 ( .B(n3591), .A(n3568), .S(n3588), .Y(n5405) );
  MUX2X1 U331 ( .B(n3592), .A(n3570), .S(n3588), .Y(n5404) );
  MUX2X1 U332 ( .B(n3593), .A(n3572), .S(n3588), .Y(n5403) );
  MUX2X1 U333 ( .B(n3594), .A(n3574), .S(n3588), .Y(n5402) );
  MUX2X1 U334 ( .B(n3595), .A(n3576), .S(n3588), .Y(n5401) );
  OAI22X1 U335 ( .A(n3596), .B(n3597), .C(n3598), .D(n3599), .Y(n3588) );
  MUX2X1 U336 ( .B(n3600), .A(n3561), .S(n3601), .Y(n5400) );
  MUX2X1 U337 ( .B(n3602), .A(n3564), .S(n3601), .Y(n5399) );
  MUX2X1 U338 ( .B(n3603), .A(n3566), .S(n3601), .Y(n5398) );
  MUX2X1 U339 ( .B(n3604), .A(n3568), .S(n3601), .Y(n5397) );
  MUX2X1 U340 ( .B(n3605), .A(n3570), .S(n3601), .Y(n5396) );
  MUX2X1 U341 ( .B(n3606), .A(n3572), .S(n3601), .Y(n5395) );
  MUX2X1 U342 ( .B(n3607), .A(n3574), .S(n3601), .Y(n5394) );
  MUX2X1 U343 ( .B(n3608), .A(n3576), .S(n3601), .Y(n5393) );
  OAI22X1 U344 ( .A(n3596), .B(n3609), .C(n3599), .D(n3610), .Y(n3601) );
  MUX2X1 U345 ( .B(n3611), .A(n3561), .S(n3612), .Y(n5392) );
  MUX2X1 U346 ( .B(n3613), .A(n3564), .S(n3612), .Y(n5391) );
  MUX2X1 U347 ( .B(n3614), .A(n3566), .S(n3612), .Y(n5390) );
  MUX2X1 U348 ( .B(n3615), .A(n3568), .S(n3612), .Y(n5389) );
  MUX2X1 U349 ( .B(n3616), .A(n3570), .S(n3612), .Y(n5388) );
  MUX2X1 U350 ( .B(n3617), .A(n3572), .S(n3612), .Y(n5387) );
  MUX2X1 U351 ( .B(n3618), .A(n3574), .S(n3612), .Y(n5386) );
  MUX2X1 U352 ( .B(n3619), .A(n3576), .S(n3612), .Y(n5385) );
  OAI22X1 U353 ( .A(n3596), .B(n3620), .C(n3598), .D(n3621), .Y(n3612) );
  MUX2X1 U354 ( .B(n3622), .A(n3561), .S(n3623), .Y(n5384) );
  MUX2X1 U355 ( .B(n3624), .A(n3564), .S(n3623), .Y(n5383) );
  MUX2X1 U356 ( .B(n3625), .A(n3566), .S(n3623), .Y(n5382) );
  MUX2X1 U357 ( .B(n3626), .A(n3568), .S(n3623), .Y(n5381) );
  MUX2X1 U358 ( .B(n3627), .A(n3570), .S(n3623), .Y(n5380) );
  MUX2X1 U359 ( .B(n3628), .A(n3572), .S(n3623), .Y(n5379) );
  MUX2X1 U360 ( .B(n3629), .A(n3574), .S(n3623), .Y(n5378) );
  MUX2X1 U361 ( .B(n3630), .A(n3576), .S(n3623), .Y(n5377) );
  OAI22X1 U362 ( .A(n3596), .B(n3631), .C(n3610), .D(n3621), .Y(n3623) );
  MUX2X1 U363 ( .B(n3632), .A(n3561), .S(n3633), .Y(n5376) );
  MUX2X1 U364 ( .B(n3634), .A(n3564), .S(n3633), .Y(n5375) );
  MUX2X1 U365 ( .B(n3635), .A(n3566), .S(n3633), .Y(n5374) );
  MUX2X1 U366 ( .B(n3636), .A(n3568), .S(n3633), .Y(n5373) );
  MUX2X1 U367 ( .B(n3637), .A(n3570), .S(n3633), .Y(n5372) );
  MUX2X1 U368 ( .B(n3638), .A(n3572), .S(n3633), .Y(n5371) );
  MUX2X1 U369 ( .B(n3639), .A(n3574), .S(n3633), .Y(n5370) );
  MUX2X1 U370 ( .B(n3640), .A(n3576), .S(n3633), .Y(n5369) );
  OAI22X1 U371 ( .A(n3596), .B(n3641), .C(n3598), .D(n3642), .Y(n3633) );
  MUX2X1 U372 ( .B(n3643), .A(n3561), .S(n3644), .Y(n5368) );
  MUX2X1 U373 ( .B(n3645), .A(n3564), .S(n3644), .Y(n5367) );
  MUX2X1 U374 ( .B(n3646), .A(n3566), .S(n3644), .Y(n5366) );
  MUX2X1 U375 ( .B(n3647), .A(n3568), .S(n3644), .Y(n5365) );
  MUX2X1 U376 ( .B(n3648), .A(n3570), .S(n3644), .Y(n5364) );
  MUX2X1 U377 ( .B(n3649), .A(n3572), .S(n3644), .Y(n5363) );
  MUX2X1 U378 ( .B(n3650), .A(n3574), .S(n3644), .Y(n5362) );
  MUX2X1 U379 ( .B(n3651), .A(n3576), .S(n3644), .Y(n5361) );
  OAI22X1 U380 ( .A(n3596), .B(n3652), .C(n3610), .D(n3642), .Y(n3644) );
  MUX2X1 U381 ( .B(n3653), .A(n3561), .S(n3654), .Y(n5360) );
  MUX2X1 U382 ( .B(n3655), .A(n3564), .S(n3654), .Y(n5359) );
  MUX2X1 U383 ( .B(n3656), .A(n3566), .S(n3654), .Y(n5358) );
  MUX2X1 U384 ( .B(n3657), .A(n3568), .S(n3654), .Y(n5357) );
  MUX2X1 U385 ( .B(n3658), .A(n3570), .S(n3654), .Y(n5356) );
  MUX2X1 U386 ( .B(n3659), .A(n3572), .S(n3654), .Y(n5355) );
  MUX2X1 U387 ( .B(n3660), .A(n3574), .S(n3654), .Y(n5354) );
  MUX2X1 U388 ( .B(n3661), .A(n3576), .S(n3654), .Y(n5353) );
  OAI21X1 U389 ( .A(n3596), .B(n3662), .C(n3663), .Y(n3654) );
  NAND3X1 U390 ( .A(n3581), .B(n3664), .C(n3665), .Y(n3663) );
  MUX2X1 U391 ( .B(n3666), .A(n3561), .S(n3667), .Y(n5352) );
  MUX2X1 U392 ( .B(n3668), .A(n3564), .S(n3667), .Y(n5351) );
  MUX2X1 U393 ( .B(n3669), .A(n3566), .S(n3667), .Y(n5350) );
  MUX2X1 U394 ( .B(n3670), .A(n3568), .S(n3667), .Y(n5349) );
  MUX2X1 U395 ( .B(n3671), .A(n3570), .S(n3667), .Y(n5348) );
  MUX2X1 U396 ( .B(n3672), .A(n3572), .S(n3667), .Y(n5347) );
  MUX2X1 U397 ( .B(n3673), .A(n3574), .S(n3667), .Y(n5346) );
  MUX2X1 U398 ( .B(n3674), .A(n3576), .S(n3667), .Y(n5345) );
  OAI22X1 U399 ( .A(n3675), .B(n3676), .C(n3677), .D(n3596), .Y(n3667) );
  NAND3X1 U400 ( .A(n3584), .B(n3586), .C(n3678), .Y(n3596) );
  MUX2X1 U401 ( .B(n3679), .A(n3561), .S(n3680), .Y(n5344) );
  MUX2X1 U402 ( .B(n3681), .A(n3564), .S(n3680), .Y(n5343) );
  MUX2X1 U403 ( .B(n3740), .A(n3566), .S(n3680), .Y(n5342) );
  MUX2X1 U404 ( .B(n3749), .A(n3568), .S(n3680), .Y(n5341) );
  MUX2X1 U405 ( .B(n3750), .A(n3570), .S(n3680), .Y(n5340) );
  MUX2X1 U406 ( .B(n3751), .A(n3572), .S(n3680), .Y(n5339) );
  MUX2X1 U407 ( .B(n3752), .A(n3574), .S(n3680), .Y(n5338) );
  MUX2X1 U408 ( .B(n3753), .A(n3576), .S(n3680), .Y(n5337) );
  OAI22X1 U409 ( .A(n3597), .B(n3754), .C(n3599), .D(n3755), .Y(n3680) );
  MUX2X1 U410 ( .B(n3756), .A(n3561), .S(n3757), .Y(n5336) );
  INVX1 U411 ( .A(N1735), .Y(n3756) );
  MUX2X1 U412 ( .B(n3758), .A(n3564), .S(n3757), .Y(n5335) );
  MUX2X1 U413 ( .B(n3759), .A(n3566), .S(n3757), .Y(n5334) );
  MUX2X1 U414 ( .B(n3760), .A(n3568), .S(n3757), .Y(n5333) );
  MUX2X1 U415 ( .B(n3761), .A(n3570), .S(n3757), .Y(n5332) );
  MUX2X1 U416 ( .B(n3762), .A(n3572), .S(n3757), .Y(n5331) );
  MUX2X1 U417 ( .B(n3763), .A(n3574), .S(n3757), .Y(n5330) );
  MUX2X1 U418 ( .B(n3764), .A(n3576), .S(n3757), .Y(n5329) );
  OAI22X1 U419 ( .A(n3609), .B(n3754), .C(n3599), .D(n3765), .Y(n3757) );
  NAND2X1 U420 ( .A(n3581), .B(n3766), .Y(n3599) );
  MUX2X1 U421 ( .B(n3767), .A(n3576), .S(n3768), .Y(n5328) );
  MUX2X1 U422 ( .B(n3769), .A(n3561), .S(n3768), .Y(n5327) );
  MUX2X1 U423 ( .B(n3770), .A(n3564), .S(n3768), .Y(n5326) );
  MUX2X1 U424 ( .B(n3771), .A(n3566), .S(n3768), .Y(n5325) );
  MUX2X1 U425 ( .B(n3772), .A(n3568), .S(n3768), .Y(n5324) );
  MUX2X1 U426 ( .B(n3773), .A(n3570), .S(n3768), .Y(n5323) );
  MUX2X1 U427 ( .B(n3774), .A(n3572), .S(n3768), .Y(n5322) );
  MUX2X1 U428 ( .B(n3775), .A(n3574), .S(n3768), .Y(n5321) );
  OAI22X1 U429 ( .A(n3620), .B(n3754), .C(n3621), .D(n3755), .Y(n3768) );
  MUX2X1 U430 ( .B(n3776), .A(n3561), .S(n3777), .Y(n5320) );
  MUX2X1 U431 ( .B(n3778), .A(n3564), .S(n3777), .Y(n5319) );
  MUX2X1 U432 ( .B(n3779), .A(n3566), .S(n3777), .Y(n5318) );
  MUX2X1 U433 ( .B(n3780), .A(n3568), .S(n3777), .Y(n5317) );
  MUX2X1 U434 ( .B(n3781), .A(n3570), .S(n3777), .Y(n5316) );
  MUX2X1 U435 ( .B(n3782), .A(n3572), .S(n3777), .Y(n5315) );
  MUX2X1 U436 ( .B(n3783), .A(n3574), .S(n3777), .Y(n5314) );
  MUX2X1 U437 ( .B(n3784), .A(n3576), .S(n3777), .Y(n5313) );
  OAI22X1 U438 ( .A(n3631), .B(n3754), .C(n3621), .D(n3765), .Y(n3777) );
  NAND2X1 U439 ( .A(n3785), .B(n3581), .Y(n3621) );
  MUX2X1 U440 ( .B(n3786), .A(n3561), .S(n3787), .Y(n5312) );
  MUX2X1 U441 ( .B(n3788), .A(n3564), .S(n3787), .Y(n5311) );
  MUX2X1 U442 ( .B(n3789), .A(n3566), .S(n3787), .Y(n5310) );
  MUX2X1 U443 ( .B(n3790), .A(n3568), .S(n3787), .Y(n5309) );
  MUX2X1 U444 ( .B(n3791), .A(n3570), .S(n3787), .Y(n5308) );
  MUX2X1 U445 ( .B(n3792), .A(n3572), .S(n3787), .Y(n5307) );
  MUX2X1 U446 ( .B(n3793), .A(n3574), .S(n3787), .Y(n5306) );
  MUX2X1 U447 ( .B(n3794), .A(n3576), .S(n3787), .Y(n5305) );
  OAI22X1 U448 ( .A(n3641), .B(n3754), .C(n3642), .D(n3755), .Y(n3787) );
  MUX2X1 U449 ( .B(n3795), .A(n3561), .S(n3796), .Y(n5304) );
  MUX2X1 U450 ( .B(n3797), .A(n3564), .S(n3796), .Y(n5303) );
  MUX2X1 U451 ( .B(n3798), .A(n3566), .S(n3796), .Y(n5302) );
  MUX2X1 U452 ( .B(n3799), .A(n3568), .S(n3796), .Y(n5301) );
  MUX2X1 U453 ( .B(n3800), .A(n3570), .S(n3796), .Y(n5300) );
  MUX2X1 U454 ( .B(n3801), .A(n3572), .S(n3796), .Y(n5299) );
  MUX2X1 U455 ( .B(n3802), .A(n3574), .S(n3796), .Y(n5298) );
  MUX2X1 U456 ( .B(n3803), .A(n3576), .S(n3796), .Y(n5297) );
  OAI22X1 U457 ( .A(n3652), .B(n3754), .C(n3642), .D(n3765), .Y(n3796) );
  NAND2X1 U458 ( .A(n3804), .B(n3581), .Y(n3642) );
  MUX2X1 U459 ( .B(n3805), .A(n3561), .S(n3806), .Y(n5296) );
  MUX2X1 U460 ( .B(n3807), .A(n3564), .S(n3806), .Y(n5295) );
  MUX2X1 U461 ( .B(n3808), .A(n3566), .S(n3806), .Y(n5294) );
  MUX2X1 U462 ( .B(n3809), .A(n3568), .S(n3806), .Y(n5293) );
  MUX2X1 U463 ( .B(n3810), .A(n3570), .S(n3806), .Y(n5292) );
  MUX2X1 U464 ( .B(n3811), .A(n3572), .S(n3806), .Y(n5291) );
  MUX2X1 U465 ( .B(n3812), .A(n3574), .S(n3806), .Y(n5290) );
  MUX2X1 U466 ( .B(n3813), .A(n3576), .S(n3806), .Y(n5289) );
  OAI21X1 U467 ( .A(n3662), .B(n3754), .C(n3814), .Y(n3806) );
  NAND3X1 U468 ( .A(n3581), .B(n3815), .C(n3816), .Y(n3814) );
  MUX2X1 U469 ( .B(n3817), .A(n3561), .S(n3818), .Y(n5288) );
  MUX2X1 U470 ( .B(n3819), .A(n3564), .S(n3818), .Y(n5287) );
  MUX2X1 U471 ( .B(n3820), .A(n3566), .S(n3818), .Y(n5286) );
  MUX2X1 U472 ( .B(n3821), .A(n3568), .S(n3818), .Y(n5285) );
  MUX2X1 U473 ( .B(n3822), .A(n3570), .S(n3818), .Y(n5284) );
  MUX2X1 U474 ( .B(n3823), .A(n3572), .S(n3818), .Y(n5283) );
  MUX2X1 U475 ( .B(n3824), .A(n3574), .S(n3818), .Y(n5282) );
  MUX2X1 U476 ( .B(n3825), .A(n3576), .S(n3818), .Y(n5281) );
  OAI22X1 U477 ( .A(n3675), .B(n3826), .C(n3677), .D(n3754), .Y(n3818) );
  NAND3X1 U478 ( .A(n3584), .B(n3585), .C(n3827), .Y(n3754) );
  MUX2X1 U479 ( .B(n3561), .A(n3828), .S(n3829), .Y(n5280) );
  MUX2X1 U480 ( .B(n3564), .A(n3830), .S(n3829), .Y(n5279) );
  MUX2X1 U481 ( .B(n3566), .A(n3831), .S(n3829), .Y(n5278) );
  MUX2X1 U482 ( .B(n3568), .A(n3832), .S(n3829), .Y(n5277) );
  MUX2X1 U483 ( .B(n3570), .A(n3833), .S(n3829), .Y(n5276) );
  MUX2X1 U484 ( .B(n3572), .A(n3834), .S(n3829), .Y(n5275) );
  MUX2X1 U485 ( .B(n3574), .A(n3835), .S(n3829), .Y(n5274) );
  MUX2X1 U486 ( .B(n3576), .A(n3836), .S(n3829), .Y(n5273) );
  AOI22X1 U487 ( .A(n3581), .B(n3837), .C(n3838), .D(n3839), .Y(n3829) );
  INVX1 U488 ( .A(n3840), .Y(n3837) );
  MUX2X1 U489 ( .B(n3841), .A(n3561), .S(n3842), .Y(n5272) );
  MUX2X1 U490 ( .B(n3843), .A(n3564), .S(n3842), .Y(n5271) );
  MUX2X1 U491 ( .B(n3844), .A(n3566), .S(n3842), .Y(n5270) );
  MUX2X1 U492 ( .B(n3845), .A(n3568), .S(n3842), .Y(n5269) );
  MUX2X1 U493 ( .B(n3846), .A(n3570), .S(n3842), .Y(n5268) );
  MUX2X1 U494 ( .B(n3847), .A(n3572), .S(n3842), .Y(n5267) );
  MUX2X1 U495 ( .B(n3848), .A(n3574), .S(n3842), .Y(n5266) );
  MUX2X1 U496 ( .B(n3849), .A(n3576), .S(n3842), .Y(n5265) );
  OAI21X1 U497 ( .A(n3850), .B(n3851), .C(n3852), .Y(n3842) );
  NAND3X1 U498 ( .A(n3853), .B(n3854), .C(n3855), .Y(n3852) );
  NOR2X1 U499 ( .A(n3856), .B(n3857), .Y(n3855) );
  INVX1 U500 ( .A(rst_b), .Y(n3856) );
  OAI21X1 U501 ( .A(n3858), .B(n3859), .C(n7246), .Y(n3851) );
  OAI21X1 U502 ( .A(n3860), .B(n3861), .C(N2777), .Y(n3859) );
  INVX1 U503 ( .A(n3853), .Y(n3861) );
  OAI21X1 U504 ( .A(n3862), .B(n3863), .C(n3864), .Y(n3858) );
  NAND2X1 U505 ( .A(n3865), .B(n3866), .Y(n3863) );
  MUX2X1 U506 ( .B(n3561), .A(n3867), .S(n3868), .Y(n5264) );
  INVX1 U507 ( .A(\regX[5][0] ), .Y(n3867) );
  MUX2X1 U508 ( .B(n3564), .A(n3869), .S(n3868), .Y(n5263) );
  INVX1 U509 ( .A(\regX[5][1] ), .Y(n3869) );
  MUX2X1 U510 ( .B(n3566), .A(n3870), .S(n3868), .Y(n5262) );
  INVX1 U511 ( .A(\regX[5][2] ), .Y(n3870) );
  MUX2X1 U512 ( .B(n3568), .A(n3871), .S(n3868), .Y(n5261) );
  INVX1 U513 ( .A(\regX[5][3] ), .Y(n3871) );
  MUX2X1 U514 ( .B(n3570), .A(n3872), .S(n3868), .Y(n5260) );
  MUX2X1 U515 ( .B(n3572), .A(n3873), .S(n3868), .Y(n5259) );
  MUX2X1 U516 ( .B(n3574), .A(n3874), .S(n3868), .Y(n5258) );
  MUX2X1 U517 ( .B(n3576), .A(n3875), .S(n3868), .Y(n5257) );
  AOI22X1 U518 ( .A(n3581), .B(n3876), .C(n3584), .D(n3877), .Y(n3868) );
  INVX1 U519 ( .A(n3878), .Y(n3584) );
  MUX2X1 U520 ( .B(n3561), .A(n3879), .S(n3880), .Y(n5256) );
  MUX2X1 U521 ( .B(n3564), .A(n3881), .S(n3880), .Y(n5255) );
  MUX2X1 U522 ( .B(n3566), .A(n3882), .S(n3880), .Y(n5254) );
  MUX2X1 U523 ( .B(n3568), .A(n3883), .S(n3880), .Y(n5253) );
  MUX2X1 U524 ( .B(n3570), .A(n3884), .S(n3880), .Y(n5252) );
  MUX2X1 U525 ( .B(n3572), .A(n3885), .S(n3880), .Y(n5251) );
  MUX2X1 U526 ( .B(n3574), .A(n3886), .S(n3880), .Y(n5250) );
  MUX2X1 U527 ( .B(n3576), .A(n3887), .S(n3880), .Y(n5249) );
  AOI22X1 U528 ( .A(n3581), .B(n3888), .C(n3889), .D(n3839), .Y(n3880) );
  INVX1 U529 ( .A(n3890), .Y(n3888) );
  MUX2X1 U530 ( .B(n3561), .A(n3891), .S(n3892), .Y(n5248) );
  MUX2X1 U531 ( .B(n3564), .A(n3893), .S(n3892), .Y(n5247) );
  MUX2X1 U532 ( .B(n3566), .A(n3894), .S(n3892), .Y(n5246) );
  MUX2X1 U533 ( .B(n3568), .A(n3895), .S(n3892), .Y(n5245) );
  MUX2X1 U534 ( .B(n3570), .A(n3896), .S(n3892), .Y(n5244) );
  MUX2X1 U535 ( .B(n3572), .A(n3897), .S(n3892), .Y(n5243) );
  MUX2X1 U536 ( .B(n3574), .A(n3898), .S(n3892), .Y(n5242) );
  MUX2X1 U537 ( .B(n3576), .A(n3899), .S(n3892), .Y(n5241) );
  AOI22X1 U538 ( .A(n3581), .B(n3900), .C(n3901), .D(n3839), .Y(n3892) );
  INVX1 U539 ( .A(n3902), .Y(n3900) );
  MUX2X1 U540 ( .B(n3903), .A(n3561), .S(n3904), .Y(n5240) );
  MUX2X1 U541 ( .B(n3905), .A(n3564), .S(n3904), .Y(n5239) );
  MUX2X1 U542 ( .B(n3906), .A(n3566), .S(n3904), .Y(n5238) );
  MUX2X1 U543 ( .B(n3907), .A(n3568), .S(n3904), .Y(n5237) );
  MUX2X1 U544 ( .B(n3908), .A(n3570), .S(n3904), .Y(n5236) );
  MUX2X1 U545 ( .B(n3909), .A(n3572), .S(n3904), .Y(n5235) );
  MUX2X1 U546 ( .B(n3910), .A(n3574), .S(n3904), .Y(n5234) );
  MUX2X1 U547 ( .B(n3911), .A(n3576), .S(n3904), .Y(n5233) );
  OAI22X1 U548 ( .A(n3675), .B(n3912), .C(n3878), .D(n3913), .Y(n3904) );
  MUX2X1 U549 ( .B(n3561), .A(n3914), .S(n3915), .Y(n5232) );
  MUX2X1 U550 ( .B(n3564), .A(n3916), .S(n3915), .Y(n5231) );
  MUX2X1 U551 ( .B(n3566), .A(n3917), .S(n3915), .Y(n5230) );
  MUX2X1 U552 ( .B(n3568), .A(n3918), .S(n3915), .Y(n5229) );
  MUX2X1 U553 ( .B(n3570), .A(n3919), .S(n3915), .Y(n5228) );
  MUX2X1 U554 ( .B(n3572), .A(n3920), .S(n3915), .Y(n5227) );
  MUX2X1 U555 ( .B(n3574), .A(n3921), .S(n3915), .Y(n5226) );
  MUX2X1 U556 ( .B(n3576), .A(n3922), .S(n3915), .Y(n5225) );
  AOI22X1 U557 ( .A(n3581), .B(n3923), .C(n3924), .D(n3839), .Y(n3915) );
  INVX1 U558 ( .A(n3925), .Y(n3923) );
  MUX2X1 U559 ( .B(n3566), .A(n3926), .S(n3927), .Y(n5224) );
  NAND2X1 U560 ( .A(InData[2]), .B(n3490), .Y(n3566) );
  MUX2X1 U561 ( .B(n3568), .A(n3928), .S(n3927), .Y(n5223) );
  NAND2X1 U562 ( .A(InData[3]), .B(n3490), .Y(n3568) );
  MUX2X1 U563 ( .B(n3570), .A(n3929), .S(n3927), .Y(n5222) );
  NAND2X1 U564 ( .A(InData[4]), .B(n3490), .Y(n3570) );
  MUX2X1 U565 ( .B(n3572), .A(n3930), .S(n3927), .Y(n5221) );
  NAND2X1 U566 ( .A(InData[5]), .B(n3490), .Y(n3572) );
  MUX2X1 U567 ( .B(n3574), .A(n3931), .S(n3927), .Y(n5220) );
  NAND2X1 U568 ( .A(InData[6]), .B(n3490), .Y(n3574) );
  MUX2X1 U569 ( .B(n3576), .A(n3932), .S(n3927), .Y(n5219) );
  NAND2X1 U570 ( .A(InData[7]), .B(n3490), .Y(n3576) );
  MUX2X1 U571 ( .B(n3561), .A(n3933), .S(n3927), .Y(n5218) );
  NAND2X1 U572 ( .A(InData[0]), .B(n3490), .Y(n3561) );
  MUX2X1 U573 ( .B(n3564), .A(n3934), .S(n3927), .Y(n5217) );
  AOI22X1 U574 ( .A(n3581), .B(n3935), .C(n3583), .D(n3839), .Y(n3927) );
  NOR2X1 U575 ( .A(n3862), .B(n3878), .Y(n3839) );
  NAND3X1 U576 ( .A(n3936), .B(n3866), .C(n7204), .Y(n3878) );
  XOR2X1 U577 ( .A(N3194), .B(n3937), .Y(n3866) );
  NOR2X1 U578 ( .A(n3938), .B(n3939), .Y(n3937) );
  INVX1 U579 ( .A(n3940), .Y(n3939) );
  INVX1 U580 ( .A(n3941), .Y(n3935) );
  INVX1 U581 ( .A(n3675), .Y(n3581) );
  NAND3X1 U582 ( .A(n3853), .B(n3942), .C(rst_b), .Y(n3675) );
  OAI21X1 U583 ( .A(n3550), .B(n3943), .C(n3857), .Y(n3942) );
  NAND3X1 U584 ( .A(n3490), .B(n3944), .C(n3945), .Y(n3857) );
  INVX1 U585 ( .A(n3545), .Y(n3550) );
  NAND2X1 U586 ( .A(InData[1]), .B(n3490), .Y(n3564) );
  OAI21X1 U587 ( .A(n3946), .B(n3947), .C(n3948), .Y(n5216) );
  NAND2X1 U588 ( .A(N2513), .B(n3949), .Y(n3948) );
  OAI21X1 U589 ( .A(n3946), .B(n3950), .C(n3951), .Y(n5215) );
  NAND2X1 U590 ( .A(N2514), .B(n3949), .Y(n3951) );
  OAI21X1 U591 ( .A(n3946), .B(n3952), .C(n3953), .Y(n5214) );
  NAND2X1 U592 ( .A(N2515), .B(n3949), .Y(n3953) );
  OAI21X1 U593 ( .A(n3946), .B(n3954), .C(n3955), .Y(n5213) );
  NAND2X1 U594 ( .A(N2516), .B(n3949), .Y(n3955) );
  OAI21X1 U595 ( .A(n3946), .B(n3956), .C(n3957), .Y(n5212) );
  NAND2X1 U596 ( .A(N2517), .B(n3949), .Y(n3957) );
  OAI21X1 U597 ( .A(n3946), .B(n3958), .C(n3959), .Y(n5211) );
  NAND2X1 U598 ( .A(N2518), .B(n3949), .Y(n3959) );
  OAI21X1 U599 ( .A(n3946), .B(n3960), .C(n3961), .Y(n5210) );
  NAND2X1 U600 ( .A(N2519), .B(n3949), .Y(n3961) );
  OAI21X1 U601 ( .A(n3946), .B(n3962), .C(n3963), .Y(n5209) );
  NAND2X1 U602 ( .A(N2520), .B(n3949), .Y(n3963) );
  OAI21X1 U603 ( .A(n3946), .B(n3964), .C(n3965), .Y(n5208) );
  NAND2X1 U604 ( .A(N2521), .B(n3949), .Y(n3965) );
  OAI21X1 U605 ( .A(n3946), .B(n3966), .C(n3967), .Y(n5207) );
  NAND2X1 U606 ( .A(N2522), .B(n3949), .Y(n3967) );
  OAI21X1 U607 ( .A(n3946), .B(n3968), .C(n3969), .Y(n5206) );
  NAND2X1 U608 ( .A(N2523), .B(n3949), .Y(n3969) );
  OAI21X1 U609 ( .A(n3946), .B(n3970), .C(n3971), .Y(n5205) );
  NAND2X1 U610 ( .A(N2524), .B(n3949), .Y(n3971) );
  INVX1 U611 ( .A(Gy[11]), .Y(n3970) );
  OAI21X1 U612 ( .A(n3946), .B(n3972), .C(n3973), .Y(n5204) );
  NAND2X1 U613 ( .A(N2525), .B(n3949), .Y(n3973) );
  INVX1 U614 ( .A(Gy[12]), .Y(n3972) );
  OAI21X1 U615 ( .A(n3946), .B(n3974), .C(n3975), .Y(n5203) );
  NAND2X1 U616 ( .A(N2526), .B(n3949), .Y(n3975) );
  INVX1 U617 ( .A(Gy[13]), .Y(n3974) );
  OAI21X1 U618 ( .A(n3946), .B(n3976), .C(n3977), .Y(n5202) );
  NAND2X1 U619 ( .A(N2527), .B(n3949), .Y(n3977) );
  INVX1 U620 ( .A(Gy[14]), .Y(n3976) );
  OAI21X1 U621 ( .A(n3946), .B(n3978), .C(n3979), .Y(n5201) );
  NAND2X1 U622 ( .A(N2528), .B(n3949), .Y(n3979) );
  INVX1 U623 ( .A(Gy[15]), .Y(n3978) );
  OAI21X1 U624 ( .A(n3946), .B(n3980), .C(n3981), .Y(n5200) );
  NAND2X1 U625 ( .A(N2529), .B(n3949), .Y(n3981) );
  INVX1 U626 ( .A(Gy[16]), .Y(n3980) );
  OAI21X1 U627 ( .A(n3946), .B(n3982), .C(n3983), .Y(n5199) );
  NAND2X1 U628 ( .A(N2530), .B(n3949), .Y(n3983) );
  INVX1 U629 ( .A(Gy[17]), .Y(n3982) );
  OAI21X1 U630 ( .A(n3946), .B(n3984), .C(n3985), .Y(n5198) );
  NAND2X1 U631 ( .A(N2531), .B(n3949), .Y(n3985) );
  INVX1 U632 ( .A(Gy[18]), .Y(n3984) );
  OAI21X1 U633 ( .A(n3946), .B(n3986), .C(n3987), .Y(n5197) );
  NAND2X1 U634 ( .A(N2532), .B(n3949), .Y(n3987) );
  INVX1 U635 ( .A(Gy[19]), .Y(n3986) );
  OAI21X1 U636 ( .A(n3946), .B(n3988), .C(n3989), .Y(n5196) );
  NAND2X1 U637 ( .A(N2533), .B(n3949), .Y(n3989) );
  INVX1 U638 ( .A(Gy[20]), .Y(n3988) );
  OAI21X1 U639 ( .A(n3946), .B(n3990), .C(n3991), .Y(n5195) );
  NAND2X1 U640 ( .A(N2534), .B(n3949), .Y(n3991) );
  INVX1 U641 ( .A(Gy[21]), .Y(n3990) );
  OAI21X1 U642 ( .A(n3946), .B(n3992), .C(n3993), .Y(n5194) );
  NAND2X1 U643 ( .A(N2535), .B(n3949), .Y(n3993) );
  INVX1 U644 ( .A(Gy[22]), .Y(n3992) );
  OAI21X1 U645 ( .A(n3946), .B(n3994), .C(n3995), .Y(n5193) );
  NAND2X1 U646 ( .A(N2536), .B(n3949), .Y(n3995) );
  INVX1 U647 ( .A(Gy[23]), .Y(n3994) );
  OAI21X1 U648 ( .A(n3946), .B(n3996), .C(n3997), .Y(n5192) );
  NAND2X1 U649 ( .A(N2537), .B(n3949), .Y(n3997) );
  INVX1 U650 ( .A(Gy[24]), .Y(n3996) );
  OAI21X1 U651 ( .A(n3946), .B(n3998), .C(n3999), .Y(n5191) );
  NAND2X1 U652 ( .A(N2538), .B(n3949), .Y(n3999) );
  INVX1 U653 ( .A(Gy[25]), .Y(n3998) );
  OAI21X1 U654 ( .A(n3946), .B(n4000), .C(n4001), .Y(n5190) );
  NAND2X1 U655 ( .A(N2539), .B(n3949), .Y(n4001) );
  INVX1 U656 ( .A(Gy[26]), .Y(n4000) );
  OAI21X1 U657 ( .A(n3946), .B(n4002), .C(n4003), .Y(n5189) );
  NAND2X1 U658 ( .A(N2540), .B(n3949), .Y(n4003) );
  INVX1 U659 ( .A(Gy[27]), .Y(n4002) );
  OAI21X1 U660 ( .A(n3946), .B(n4004), .C(n4005), .Y(n5188) );
  NAND2X1 U661 ( .A(N2541), .B(n3949), .Y(n4005) );
  INVX1 U662 ( .A(Gy[28]), .Y(n4004) );
  OAI21X1 U663 ( .A(n3946), .B(n4006), .C(n4007), .Y(n5187) );
  NAND2X1 U664 ( .A(N2542), .B(n3949), .Y(n4007) );
  INVX1 U665 ( .A(Gy[29]), .Y(n4006) );
  OAI21X1 U666 ( .A(n3946), .B(n4008), .C(n4009), .Y(n5186) );
  NAND2X1 U667 ( .A(N2543), .B(n3949), .Y(n4009) );
  INVX1 U668 ( .A(Gy[30]), .Y(n4008) );
  OAI21X1 U669 ( .A(n3946), .B(n4010), .C(n4011), .Y(n5185) );
  NAND2X1 U670 ( .A(N2544), .B(n3949), .Y(n4011) );
  INVX1 U671 ( .A(n4012), .Y(n3949) );
  INVX1 U672 ( .A(Gy[31]), .Y(n4010) );
  OAI21X1 U673 ( .A(n7282), .B(n3555), .C(n4013), .Y(n5152) );
  AOI22X1 U674 ( .A(N2300), .B(n4014), .C(Gx[0]), .D(n4015), .Y(n4013) );
  INVX1 U675 ( .A(N4393), .Y(n7282) );
  OAI21X1 U676 ( .A(n7291), .B(n3555), .C(n4016), .Y(n5151) );
  AOI22X1 U677 ( .A(N2301), .B(n4014), .C(Gx[1]), .D(n4015), .Y(n4016) );
  INVX1 U678 ( .A(N4390), .Y(n7291) );
  OAI21X1 U679 ( .A(n7292), .B(n3555), .C(n4017), .Y(n5150) );
  AOI22X1 U680 ( .A(N2302), .B(n4014), .C(Gx[2]), .D(n4015), .Y(n4017) );
  INVX1 U681 ( .A(N4387), .Y(n7292) );
  OAI21X1 U682 ( .A(n7293), .B(n3555), .C(n4018), .Y(n5149) );
  AOI22X1 U683 ( .A(N2303), .B(n4014), .C(Gx[3]), .D(n4015), .Y(n4018) );
  INVX1 U684 ( .A(N4384), .Y(n7293) );
  OAI21X1 U685 ( .A(n7294), .B(n3555), .C(n4019), .Y(n5148) );
  AOI22X1 U686 ( .A(N2304), .B(n4014), .C(Gx[4]), .D(n4015), .Y(n4019) );
  INVX1 U687 ( .A(N4381), .Y(n7294) );
  OAI21X1 U688 ( .A(n7295), .B(n3555), .C(n4020), .Y(n5147) );
  AOI22X1 U689 ( .A(N2305), .B(n4014), .C(Gx[5]), .D(n4015), .Y(n4020) );
  INVX1 U690 ( .A(N4378), .Y(n7295) );
  OAI21X1 U691 ( .A(n7296), .B(n3555), .C(n4021), .Y(n5146) );
  AOI22X1 U692 ( .A(N2306), .B(n4014), .C(Gx[6]), .D(n4015), .Y(n4021) );
  INVX1 U693 ( .A(N4375), .Y(n7296) );
  OAI21X1 U694 ( .A(n7297), .B(n3555), .C(n4022), .Y(n5145) );
  AOI22X1 U695 ( .A(N2307), .B(n4014), .C(Gx[7]), .D(n4015), .Y(n4022) );
  INVX1 U696 ( .A(N4372), .Y(n7297) );
  OAI21X1 U697 ( .A(n3555), .B(n4023), .C(n4024), .Y(n5144) );
  AOI22X1 U698 ( .A(N2308), .B(n3472), .C(Gx[8]), .D(n4025), .Y(n4024) );
  OAI21X1 U699 ( .A(n3555), .B(n4026), .C(n4027), .Y(n5143) );
  AOI22X1 U700 ( .A(N2309), .B(n3472), .C(Gx[9]), .D(n4025), .Y(n4027) );
  OAI21X1 U701 ( .A(n3555), .B(n4028), .C(n4029), .Y(n5142) );
  AOI22X1 U702 ( .A(N2310), .B(n3472), .C(Gx[10]), .D(n4025), .Y(n4029) );
  OAI21X1 U703 ( .A(n3555), .B(n4030), .C(n4031), .Y(n5141) );
  AOI22X1 U704 ( .A(N2311), .B(n3472), .C(Gx[11]), .D(n4025), .Y(n4031) );
  OAI21X1 U705 ( .A(n3555), .B(n4032), .C(n4033), .Y(n5140) );
  AOI22X1 U706 ( .A(N2312), .B(n3472), .C(Gx[12]), .D(n4025), .Y(n4033) );
  OAI21X1 U707 ( .A(n3555), .B(n4034), .C(n4035), .Y(n5139) );
  AOI22X1 U708 ( .A(N2313), .B(n3472), .C(Gx[13]), .D(n4025), .Y(n4035) );
  OAI21X1 U709 ( .A(n3555), .B(n4036), .C(n4037), .Y(n5138) );
  AOI22X1 U710 ( .A(N2314), .B(n3472), .C(Gx[14]), .D(n4025), .Y(n4037) );
  OAI21X1 U711 ( .A(n3555), .B(n4038), .C(n4039), .Y(n5137) );
  AOI22X1 U712 ( .A(N2315), .B(n3472), .C(Gx[15]), .D(n4025), .Y(n4039) );
  OAI21X1 U713 ( .A(n3555), .B(n4040), .C(n4041), .Y(n5136) );
  AOI22X1 U714 ( .A(N2316), .B(n3472), .C(Gx[16]), .D(n4025), .Y(n4041) );
  OAI21X1 U715 ( .A(n3555), .B(n4042), .C(n4043), .Y(n5135) );
  AOI22X1 U716 ( .A(N2317), .B(n3472), .C(Gx[17]), .D(n4025), .Y(n4043) );
  OAI21X1 U717 ( .A(n3555), .B(n4044), .C(n4045), .Y(n5134) );
  AOI22X1 U718 ( .A(N2318), .B(n3472), .C(Gx[18]), .D(n4025), .Y(n4045) );
  OAI21X1 U719 ( .A(n3555), .B(n4046), .C(n4047), .Y(n5133) );
  AOI22X1 U720 ( .A(N2319), .B(n3472), .C(Gx[19]), .D(n4025), .Y(n4047) );
  OAI21X1 U721 ( .A(n3555), .B(n4048), .C(n4049), .Y(n5132) );
  AOI22X1 U722 ( .A(N2320), .B(n3472), .C(Gx[20]), .D(n4025), .Y(n4049) );
  OAI21X1 U723 ( .A(n3555), .B(n4050), .C(n4051), .Y(n5131) );
  AOI22X1 U724 ( .A(N2321), .B(n3472), .C(Gx[21]), .D(n4025), .Y(n4051) );
  OAI21X1 U725 ( .A(n3555), .B(n4052), .C(n4053), .Y(n5130) );
  AOI22X1 U726 ( .A(N2322), .B(n3472), .C(Gx[22]), .D(n4025), .Y(n4053) );
  OAI21X1 U727 ( .A(n3555), .B(n4054), .C(n4055), .Y(n5129) );
  AOI22X1 U728 ( .A(N2323), .B(n3472), .C(Gx[23]), .D(n4025), .Y(n4055) );
  OAI21X1 U729 ( .A(n3555), .B(n4056), .C(n4057), .Y(n5128) );
  AOI22X1 U730 ( .A(N2324), .B(n3472), .C(Gx[24]), .D(n4025), .Y(n4057) );
  OAI21X1 U731 ( .A(n3555), .B(n4058), .C(n4059), .Y(n5127) );
  AOI22X1 U732 ( .A(N2325), .B(n3472), .C(Gx[25]), .D(n4025), .Y(n4059) );
  OAI21X1 U733 ( .A(n3555), .B(n4060), .C(n4061), .Y(n5126) );
  AOI22X1 U734 ( .A(N2326), .B(n3472), .C(Gx[26]), .D(n4025), .Y(n4061) );
  OAI21X1 U735 ( .A(n3555), .B(n4062), .C(n4063), .Y(n5125) );
  AOI22X1 U736 ( .A(N2327), .B(n3472), .C(Gx[27]), .D(n4025), .Y(n4063) );
  OAI21X1 U737 ( .A(n3555), .B(n4064), .C(n4065), .Y(n5124) );
  AOI22X1 U738 ( .A(N2328), .B(n3472), .C(Gx[28]), .D(n4025), .Y(n4065) );
  OAI21X1 U739 ( .A(n3555), .B(n4066), .C(n4067), .Y(n5123) );
  AOI22X1 U740 ( .A(N2329), .B(n3472), .C(Gx[29]), .D(n4025), .Y(n4067) );
  OAI21X1 U741 ( .A(n3555), .B(n4068), .C(n4069), .Y(n5122) );
  AOI22X1 U742 ( .A(N2330), .B(n3472), .C(Gx[30]), .D(n4025), .Y(n4069) );
  OAI21X1 U743 ( .A(n3555), .B(n4070), .C(n4071), .Y(n5121) );
  AOI22X1 U744 ( .A(N2331), .B(n3472), .C(Gx[31]), .D(n4025), .Y(n4071) );
  OAI21X1 U745 ( .A(n7283), .B(n3555), .C(n4072), .Y(n5120) );
  AOI22X1 U746 ( .A(N2648), .B(n4014), .C(n4015), .D(Gy[0]), .Y(n4072) );
  INVX1 U747 ( .A(N4465), .Y(n7283) );
  OAI21X1 U748 ( .A(n7284), .B(n3555), .C(n4073), .Y(n5119) );
  AOI22X1 U749 ( .A(N2746), .B(n4014), .C(n4015), .D(Gy[1]), .Y(n4073) );
  INVX1 U750 ( .A(N4462), .Y(n7284) );
  OAI21X1 U751 ( .A(n7285), .B(n3555), .C(n4074), .Y(n5118) );
  AOI22X1 U752 ( .A(N2747), .B(n4014), .C(n4015), .D(Gy[2]), .Y(n4074) );
  INVX1 U753 ( .A(N4459), .Y(n7285) );
  OAI21X1 U754 ( .A(n7286), .B(n3555), .C(n4075), .Y(n5117) );
  AOI22X1 U755 ( .A(N2748), .B(n4014), .C(n4015), .D(Gy[3]), .Y(n4075) );
  INVX1 U756 ( .A(N4456), .Y(n7286) );
  OAI21X1 U757 ( .A(n7287), .B(n3555), .C(n4076), .Y(n5116) );
  AOI22X1 U758 ( .A(N2749), .B(n4014), .C(n4015), .D(Gy[4]), .Y(n4076) );
  INVX1 U759 ( .A(N4453), .Y(n7287) );
  OAI21X1 U760 ( .A(n7288), .B(n3555), .C(n4077), .Y(n5115) );
  AOI22X1 U761 ( .A(n4014), .B(N2750), .C(n4015), .D(Gy[5]), .Y(n4077) );
  INVX1 U762 ( .A(N4450), .Y(n7288) );
  OAI21X1 U763 ( .A(n7289), .B(n3555), .C(n4078), .Y(n5114) );
  AOI22X1 U764 ( .A(n4014), .B(N2751), .C(n4015), .D(Gy[6]), .Y(n4078) );
  INVX1 U765 ( .A(N4447), .Y(n7289) );
  OAI21X1 U766 ( .A(n7290), .B(n3555), .C(n4079), .Y(n5113) );
  AOI22X1 U767 ( .A(n4014), .B(N2752), .C(n4015), .D(Gy[7]), .Y(n4079) );
  NOR2X1 U768 ( .A(n3488), .B(n4080), .Y(n4014) );
  INVX1 U769 ( .A(N4444), .Y(n7290) );
  OAI21X1 U770 ( .A(n3555), .B(n4081), .C(n4082), .Y(n5112) );
  AOI22X1 U771 ( .A(N2753), .B(n3472), .C(n4025), .D(Gy[8]), .Y(n4082) );
  OAI21X1 U772 ( .A(n3555), .B(n4083), .C(n4084), .Y(n5111) );
  AOI22X1 U773 ( .A(N2754), .B(n3472), .C(n4025), .D(Gy[9]), .Y(n4084) );
  OAI21X1 U774 ( .A(n3555), .B(n4085), .C(n4086), .Y(n5110) );
  AOI22X1 U775 ( .A(N2755), .B(n3472), .C(n4025), .D(Gy[10]), .Y(n4086) );
  OAI21X1 U776 ( .A(n3555), .B(n4087), .C(n4088), .Y(n5109) );
  AOI22X1 U777 ( .A(N2756), .B(n3472), .C(n4025), .D(Gy[11]), .Y(n4088) );
  OAI21X1 U778 ( .A(n3555), .B(n4089), .C(n4090), .Y(n5108) );
  AOI22X1 U779 ( .A(N2757), .B(n3472), .C(n4025), .D(Gy[12]), .Y(n4090) );
  OAI21X1 U780 ( .A(n3555), .B(n4091), .C(n4092), .Y(n5107) );
  AOI22X1 U781 ( .A(N2758), .B(n3472), .C(n4025), .D(Gy[13]), .Y(n4092) );
  OAI21X1 U782 ( .A(n3555), .B(n4093), .C(n4094), .Y(n5106) );
  AOI22X1 U783 ( .A(N2759), .B(n3472), .C(n4025), .D(Gy[14]), .Y(n4094) );
  OAI21X1 U784 ( .A(n3555), .B(n4095), .C(n4096), .Y(n5105) );
  AOI22X1 U785 ( .A(N2760), .B(n3472), .C(n4025), .D(Gy[15]), .Y(n4096) );
  OAI21X1 U786 ( .A(n3555), .B(n4097), .C(n4098), .Y(n5104) );
  AOI22X1 U787 ( .A(N2761), .B(n3472), .C(n4025), .D(Gy[16]), .Y(n4098) );
  OAI21X1 U788 ( .A(n3555), .B(n4099), .C(n4100), .Y(n5103) );
  AOI22X1 U789 ( .A(N2762), .B(n3472), .C(n4025), .D(Gy[17]), .Y(n4100) );
  OAI21X1 U790 ( .A(n3555), .B(n4101), .C(n4102), .Y(n5102) );
  AOI22X1 U791 ( .A(N2763), .B(n3472), .C(n4025), .D(Gy[18]), .Y(n4102) );
  OAI21X1 U792 ( .A(n3555), .B(n4103), .C(n4104), .Y(n5101) );
  AOI22X1 U793 ( .A(N2764), .B(n3472), .C(n4025), .D(Gy[19]), .Y(n4104) );
  OAI21X1 U794 ( .A(n3555), .B(n4105), .C(n4106), .Y(n5100) );
  AOI22X1 U795 ( .A(N2765), .B(n3472), .C(n4025), .D(Gy[20]), .Y(n4106) );
  OAI21X1 U796 ( .A(n3555), .B(n4107), .C(n4108), .Y(n5099) );
  AOI22X1 U797 ( .A(N2766), .B(n3472), .C(n4025), .D(Gy[21]), .Y(n4108) );
  OAI21X1 U798 ( .A(n3555), .B(n4109), .C(n4110), .Y(n5098) );
  AOI22X1 U799 ( .A(N2767), .B(n3472), .C(n4025), .D(Gy[22]), .Y(n4110) );
  OAI21X1 U800 ( .A(n3555), .B(n4111), .C(n4112), .Y(n5097) );
  AOI22X1 U801 ( .A(N2768), .B(n3472), .C(n4025), .D(Gy[23]), .Y(n4112) );
  OAI21X1 U802 ( .A(n3555), .B(n4113), .C(n4114), .Y(n5096) );
  AOI22X1 U803 ( .A(N2769), .B(n3472), .C(n4025), .D(Gy[24]), .Y(n4114) );
  OAI21X1 U804 ( .A(n3555), .B(n4115), .C(n4116), .Y(n5095) );
  AOI22X1 U805 ( .A(N2770), .B(n3472), .C(n4025), .D(Gy[25]), .Y(n4116) );
  OAI21X1 U806 ( .A(n3555), .B(n4117), .C(n4118), .Y(n5094) );
  AOI22X1 U807 ( .A(N2771), .B(n3472), .C(n4025), .D(Gy[26]), .Y(n4118) );
  OAI21X1 U808 ( .A(n3555), .B(n4119), .C(n4120), .Y(n5093) );
  AOI22X1 U809 ( .A(N2772), .B(n3472), .C(n4025), .D(Gy[27]), .Y(n4120) );
  OAI21X1 U810 ( .A(n3555), .B(n4121), .C(n4122), .Y(n5092) );
  AOI22X1 U811 ( .A(N2773), .B(n3472), .C(n4025), .D(Gy[28]), .Y(n4122) );
  OAI21X1 U812 ( .A(n3555), .B(n4123), .C(n4124), .Y(n5091) );
  AOI22X1 U813 ( .A(N2774), .B(n3472), .C(n4025), .D(Gy[29]), .Y(n4124) );
  OAI21X1 U814 ( .A(n3555), .B(n4125), .C(n4126), .Y(n5090) );
  AOI22X1 U815 ( .A(N2775), .B(n3472), .C(n4025), .D(Gy[30]), .Y(n4126) );
  NOR2X1 U816 ( .A(n4128), .B(n3488), .Y(n4015) );
  OAI21X1 U817 ( .A(n3557), .B(n4129), .C(rst_b), .Y(n3488) );
  NOR2X1 U818 ( .A(n3547), .B(n4130), .Y(n4129) );
  NAND2X1 U819 ( .A(n3545), .B(n4131), .Y(n4130) );
  MUX2X1 U820 ( .B(n7529), .A(n4132), .S(n4133), .Y(n5088) );
  INVX1 U821 ( .A(N4369), .Y(n7529) );
  MUX2X1 U822 ( .B(n7528), .A(n4134), .S(n4133), .Y(n5087) );
  INVX1 U823 ( .A(N4366), .Y(n7528) );
  MUX2X1 U824 ( .B(n7527), .A(n4135), .S(n4133), .Y(n5086) );
  INVX1 U825 ( .A(N4363), .Y(n7527) );
  MUX2X1 U826 ( .B(n7526), .A(n4136), .S(n4133), .Y(n5085) );
  INVX1 U827 ( .A(N4360), .Y(n7526) );
  MUX2X1 U828 ( .B(n7525), .A(n4137), .S(n4133), .Y(n5084) );
  INVX1 U829 ( .A(N4357), .Y(n7525) );
  MUX2X1 U830 ( .B(n7524), .A(n4138), .S(n4133), .Y(n5083) );
  INVX1 U831 ( .A(N4354), .Y(n7524) );
  MUX2X1 U832 ( .B(n7523), .A(n4139), .S(n4133), .Y(n5082) );
  INVX1 U833 ( .A(N4351), .Y(n7523) );
  MUX2X1 U834 ( .B(n7522), .A(n4140), .S(n4133), .Y(n5081) );
  INVX1 U835 ( .A(N4348), .Y(n7522) );
  MUX2X1 U836 ( .B(n7506), .A(n4132), .S(n4141), .Y(n5080) );
  INVX1 U837 ( .A(N4345), .Y(n7506) );
  MUX2X1 U838 ( .B(n7507), .A(n4134), .S(n4141), .Y(n5079) );
  INVX1 U839 ( .A(N4342), .Y(n7507) );
  MUX2X1 U840 ( .B(n7508), .A(n4135), .S(n4141), .Y(n5078) );
  INVX1 U841 ( .A(N4339), .Y(n7508) );
  MUX2X1 U842 ( .B(n7509), .A(n4136), .S(n4141), .Y(n5077) );
  INVX1 U843 ( .A(N4336), .Y(n7509) );
  MUX2X1 U844 ( .B(n7510), .A(n4137), .S(n4141), .Y(n5076) );
  INVX1 U845 ( .A(N4333), .Y(n7510) );
  MUX2X1 U846 ( .B(n7511), .A(n4138), .S(n4141), .Y(n5075) );
  INVX1 U847 ( .A(N4330), .Y(n7511) );
  MUX2X1 U848 ( .B(n7512), .A(n4139), .S(n4141), .Y(n5074) );
  INVX1 U849 ( .A(N4327), .Y(n7512) );
  MUX2X1 U850 ( .B(n7513), .A(n4140), .S(n4141), .Y(n5073) );
  INVX1 U851 ( .A(N4324), .Y(n7513) );
  MUX2X1 U852 ( .B(n7490), .A(n4132), .S(n4142), .Y(n5072) );
  INVX1 U853 ( .A(N4321), .Y(n7490) );
  MUX2X1 U854 ( .B(n7491), .A(n4134), .S(n4142), .Y(n5071) );
  INVX1 U855 ( .A(N4318), .Y(n7491) );
  MUX2X1 U856 ( .B(n7492), .A(n4135), .S(n4142), .Y(n5070) );
  INVX1 U857 ( .A(N4315), .Y(n7492) );
  MUX2X1 U858 ( .B(n7493), .A(n4136), .S(n4142), .Y(n5069) );
  INVX1 U859 ( .A(N4312), .Y(n7493) );
  MUX2X1 U860 ( .B(n7494), .A(n4137), .S(n4142), .Y(n5068) );
  INVX1 U861 ( .A(N4309), .Y(n7494) );
  MUX2X1 U862 ( .B(n7495), .A(n4138), .S(n4142), .Y(n5067) );
  INVX1 U863 ( .A(N4306), .Y(n7495) );
  MUX2X1 U864 ( .B(n7496), .A(n4139), .S(n4142), .Y(n5066) );
  INVX1 U865 ( .A(N4303), .Y(n7496) );
  MUX2X1 U866 ( .B(n7497), .A(n4140), .S(n4142), .Y(n5065) );
  INVX1 U867 ( .A(N4300), .Y(n7497) );
  MUX2X1 U868 ( .B(n7442), .A(n4132), .S(n4143), .Y(n5064) );
  INVX1 U869 ( .A(N4297), .Y(n7442) );
  MUX2X1 U870 ( .B(n7443), .A(n4134), .S(n4143), .Y(n5063) );
  INVX1 U871 ( .A(N4294), .Y(n7443) );
  MUX2X1 U872 ( .B(n7444), .A(n4135), .S(n4143), .Y(n5062) );
  INVX1 U873 ( .A(N4291), .Y(n7444) );
  MUX2X1 U874 ( .B(n7445), .A(n4136), .S(n4143), .Y(n5061) );
  INVX1 U875 ( .A(N4288), .Y(n7445) );
  MUX2X1 U876 ( .B(n7446), .A(n4137), .S(n4143), .Y(n5060) );
  INVX1 U877 ( .A(N4285), .Y(n7446) );
  MUX2X1 U878 ( .B(n7447), .A(n4138), .S(n4143), .Y(n5059) );
  INVX1 U879 ( .A(N4282), .Y(n7447) );
  MUX2X1 U880 ( .B(n7448), .A(n4139), .S(n4143), .Y(n5058) );
  INVX1 U881 ( .A(N4279), .Y(n7448) );
  MUX2X1 U882 ( .B(n7449), .A(n4140), .S(n4143), .Y(n5057) );
  INVX1 U883 ( .A(N4276), .Y(n7449) );
  MUX2X1 U884 ( .B(n7426), .A(n4132), .S(n4144), .Y(n5056) );
  INVX1 U885 ( .A(N4273), .Y(n7426) );
  MUX2X1 U886 ( .B(n7427), .A(n4134), .S(n4144), .Y(n5055) );
  INVX1 U887 ( .A(N4270), .Y(n7427) );
  MUX2X1 U888 ( .B(n7428), .A(n4135), .S(n4144), .Y(n5054) );
  INVX1 U889 ( .A(N4267), .Y(n7428) );
  MUX2X1 U890 ( .B(n7429), .A(n4136), .S(n4144), .Y(n5053) );
  INVX1 U891 ( .A(N4264), .Y(n7429) );
  MUX2X1 U892 ( .B(n7430), .A(n4137), .S(n4144), .Y(n5052) );
  INVX1 U893 ( .A(N4261), .Y(n7430) );
  MUX2X1 U894 ( .B(n7431), .A(n4138), .S(n4144), .Y(n5051) );
  INVX1 U895 ( .A(N4258), .Y(n7431) );
  MUX2X1 U896 ( .B(n7432), .A(n4139), .S(n4144), .Y(n5050) );
  INVX1 U897 ( .A(N4255), .Y(n7432) );
  MUX2X1 U898 ( .B(n7433), .A(n4140), .S(n4144), .Y(n5049) );
  INVX1 U899 ( .A(N4252), .Y(n7433) );
  MUX2X1 U900 ( .B(n7378), .A(n4132), .S(n4145), .Y(n5048) );
  INVX1 U901 ( .A(N4249), .Y(n7378) );
  MUX2X1 U902 ( .B(n7379), .A(n4134), .S(n4145), .Y(n5047) );
  INVX1 U903 ( .A(N4246), .Y(n7379) );
  MUX2X1 U904 ( .B(n7380), .A(n4135), .S(n4145), .Y(n5046) );
  INVX1 U905 ( .A(N4243), .Y(n7380) );
  MUX2X1 U906 ( .B(n7381), .A(n4136), .S(n4145), .Y(n5045) );
  INVX1 U907 ( .A(N4240), .Y(n7381) );
  MUX2X1 U908 ( .B(n7382), .A(n4137), .S(n4145), .Y(n5044) );
  INVX1 U909 ( .A(N4237), .Y(n7382) );
  MUX2X1 U910 ( .B(n7383), .A(n4138), .S(n4145), .Y(n5043) );
  INVX1 U911 ( .A(N4234), .Y(n7383) );
  MUX2X1 U912 ( .B(n7384), .A(n4139), .S(n4145), .Y(n5042) );
  INVX1 U913 ( .A(N4231), .Y(n7384) );
  MUX2X1 U914 ( .B(n7385), .A(n4140), .S(n4145), .Y(n5041) );
  INVX1 U915 ( .A(N4228), .Y(n7385) );
  MUX2X1 U916 ( .B(n7362), .A(n4132), .S(n4146), .Y(n5040) );
  INVX1 U917 ( .A(N4225), .Y(n7362) );
  MUX2X1 U918 ( .B(n7363), .A(n4134), .S(n4146), .Y(n5039) );
  INVX1 U919 ( .A(N4222), .Y(n7363) );
  MUX2X1 U920 ( .B(n7364), .A(n4135), .S(n4146), .Y(n5038) );
  INVX1 U921 ( .A(N4219), .Y(n7364) );
  MUX2X1 U922 ( .B(n7365), .A(n4136), .S(n4146), .Y(n5037) );
  INVX1 U923 ( .A(N4216), .Y(n7365) );
  MUX2X1 U924 ( .B(n7366), .A(n4137), .S(n4146), .Y(n5036) );
  INVX1 U925 ( .A(N4213), .Y(n7366) );
  MUX2X1 U926 ( .B(n7367), .A(n4138), .S(n4146), .Y(n5035) );
  INVX1 U927 ( .A(N4210), .Y(n7367) );
  MUX2X1 U928 ( .B(n7368), .A(n4139), .S(n4146), .Y(n5034) );
  INVX1 U929 ( .A(N4207), .Y(n7368) );
  MUX2X1 U930 ( .B(n7369), .A(n4140), .S(n4146), .Y(n5033) );
  INVX1 U931 ( .A(N4204), .Y(n7369) );
  MUX2X1 U932 ( .B(n7545), .A(n4132), .S(n4147), .Y(n5032) );
  INVX1 U933 ( .A(N4201), .Y(n7545) );
  MUX2X1 U934 ( .B(n7544), .A(n4134), .S(n4147), .Y(n5031) );
  INVX1 U935 ( .A(N4198), .Y(n7544) );
  MUX2X1 U936 ( .B(n7543), .A(n4135), .S(n4147), .Y(n5030) );
  INVX1 U937 ( .A(N4195), .Y(n7543) );
  MUX2X1 U938 ( .B(n7542), .A(n4136), .S(n4147), .Y(n5029) );
  INVX1 U939 ( .A(N4192), .Y(n7542) );
  MUX2X1 U940 ( .B(n7541), .A(n4137), .S(n4147), .Y(n5028) );
  INVX1 U941 ( .A(N4189), .Y(n7541) );
  MUX2X1 U942 ( .B(n7540), .A(n4138), .S(n4147), .Y(n5027) );
  INVX1 U943 ( .A(N4186), .Y(n7540) );
  MUX2X1 U944 ( .B(n7539), .A(n4139), .S(n4147), .Y(n5026) );
  INVX1 U945 ( .A(N4183), .Y(n7539) );
  MUX2X1 U946 ( .B(n7538), .A(n4140), .S(n4147), .Y(n5025) );
  INVX1 U947 ( .A(N4180), .Y(n7538) );
  MUX2X1 U948 ( .B(n7561), .A(n4132), .S(n4148), .Y(n5024) );
  INVX1 U949 ( .A(N4177), .Y(n7561) );
  MUX2X1 U950 ( .B(n7560), .A(n4134), .S(n4148), .Y(n5023) );
  INVX1 U951 ( .A(N4174), .Y(n7560) );
  MUX2X1 U952 ( .B(n7559), .A(n4135), .S(n4148), .Y(n5022) );
  INVX1 U953 ( .A(N4171), .Y(n7559) );
  MUX2X1 U954 ( .B(n7558), .A(n4136), .S(n4148), .Y(n5021) );
  INVX1 U955 ( .A(N4168), .Y(n7558) );
  MUX2X1 U956 ( .B(n7557), .A(n4137), .S(n4148), .Y(n5020) );
  INVX1 U957 ( .A(N4165), .Y(n7557) );
  MUX2X1 U958 ( .B(n7556), .A(n4138), .S(n4148), .Y(n5019) );
  INVX1 U959 ( .A(N4162), .Y(n7556) );
  MUX2X1 U960 ( .B(n7555), .A(n4139), .S(n4148), .Y(n5018) );
  INVX1 U961 ( .A(N4159), .Y(n7555) );
  MUX2X1 U962 ( .B(n7554), .A(n4140), .S(n4148), .Y(n5017) );
  INVX1 U963 ( .A(N4156), .Y(n7554) );
  MUX2X1 U964 ( .B(n7474), .A(n4132), .S(n4149), .Y(n5016) );
  INVX1 U965 ( .A(N4153), .Y(n7474) );
  MUX2X1 U966 ( .B(n7475), .A(n4134), .S(n4149), .Y(n5015) );
  INVX1 U967 ( .A(N4150), .Y(n7475) );
  MUX2X1 U968 ( .B(n7476), .A(n4135), .S(n4149), .Y(n5014) );
  INVX1 U969 ( .A(N4147), .Y(n7476) );
  MUX2X1 U970 ( .B(n7477), .A(n4136), .S(n4149), .Y(n5013) );
  INVX1 U971 ( .A(N4144), .Y(n7477) );
  MUX2X1 U972 ( .B(n7478), .A(n4137), .S(n4149), .Y(n5012) );
  INVX1 U973 ( .A(N4141), .Y(n7478) );
  MUX2X1 U974 ( .B(n7479), .A(n4138), .S(n4149), .Y(n5011) );
  INVX1 U975 ( .A(N4138), .Y(n7479) );
  MUX2X1 U976 ( .B(n7480), .A(n4139), .S(n4149), .Y(n5010) );
  INVX1 U977 ( .A(N4135), .Y(n7480) );
  MUX2X1 U978 ( .B(n7481), .A(n4140), .S(n4149), .Y(n5009) );
  INVX1 U979 ( .A(N4132), .Y(n7481) );
  MUX2X1 U980 ( .B(n7458), .A(n4132), .S(n4150), .Y(n5008) );
  INVX1 U981 ( .A(N4129), .Y(n7458) );
  MUX2X1 U982 ( .B(n7459), .A(n4134), .S(n4150), .Y(n5007) );
  INVX1 U983 ( .A(N4126), .Y(n7459) );
  MUX2X1 U984 ( .B(n7460), .A(n4135), .S(n4150), .Y(n5006) );
  INVX1 U985 ( .A(N4123), .Y(n7460) );
  MUX2X1 U986 ( .B(n7461), .A(n4136), .S(n4150), .Y(n5005) );
  INVX1 U987 ( .A(N4120), .Y(n7461) );
  MUX2X1 U988 ( .B(n7462), .A(n4137), .S(n4150), .Y(n5004) );
  INVX1 U989 ( .A(N4117), .Y(n7462) );
  MUX2X1 U990 ( .B(n7463), .A(n4138), .S(n4150), .Y(n5003) );
  INVX1 U991 ( .A(N4114), .Y(n7463) );
  MUX2X1 U992 ( .B(n7464), .A(n4139), .S(n4150), .Y(n5002) );
  INVX1 U993 ( .A(N4111), .Y(n7464) );
  MUX2X1 U994 ( .B(n7465), .A(n4140), .S(n4150), .Y(n5001) );
  INVX1 U995 ( .A(N4108), .Y(n7465) );
  MUX2X1 U996 ( .B(n7410), .A(n4132), .S(n4151), .Y(n5000) );
  INVX1 U997 ( .A(N4105), .Y(n7410) );
  MUX2X1 U998 ( .B(n7411), .A(n4134), .S(n4151), .Y(n4999) );
  INVX1 U999 ( .A(N4102), .Y(n7411) );
  MUX2X1 U1000 ( .B(n7412), .A(n4135), .S(n4151), .Y(n4998) );
  INVX1 U1001 ( .A(N4099), .Y(n7412) );
  MUX2X1 U1002 ( .B(n7413), .A(n4136), .S(n4151), .Y(n4997) );
  INVX1 U1003 ( .A(N4096), .Y(n7413) );
  MUX2X1 U1004 ( .B(n7414), .A(n4137), .S(n4151), .Y(n4996) );
  INVX1 U1005 ( .A(N4093), .Y(n7414) );
  MUX2X1 U1006 ( .B(n7415), .A(n4138), .S(n4151), .Y(n4995) );
  INVX1 U1007 ( .A(N4090), .Y(n7415) );
  MUX2X1 U1008 ( .B(n7416), .A(n4139), .S(n4151), .Y(n4994) );
  INVX1 U1009 ( .A(N4087), .Y(n7416) );
  MUX2X1 U1010 ( .B(n7417), .A(n4140), .S(n4151), .Y(n4993) );
  INVX1 U1011 ( .A(N4084), .Y(n7417) );
  MUX2X1 U1012 ( .B(n7401), .A(n4134), .S(n4152), .Y(n4992) );
  INVX1 U1013 ( .A(N4078), .Y(n7401) );
  MUX2X1 U1014 ( .B(n7400), .A(n4135), .S(n4152), .Y(n4991) );
  INVX1 U1015 ( .A(N4075), .Y(n7400) );
  MUX2X1 U1016 ( .B(n7399), .A(n4136), .S(n4152), .Y(n4990) );
  INVX1 U1017 ( .A(N4072), .Y(n7399) );
  MUX2X1 U1018 ( .B(n7398), .A(n4137), .S(n4152), .Y(n4989) );
  INVX1 U1019 ( .A(N4069), .Y(n7398) );
  MUX2X1 U1020 ( .B(n7397), .A(n4138), .S(n4152), .Y(n4988) );
  INVX1 U1021 ( .A(N4066), .Y(n7397) );
  MUX2X1 U1022 ( .B(n7396), .A(n4139), .S(n4152), .Y(n4987) );
  INVX1 U1023 ( .A(N4063), .Y(n7396) );
  MUX2X1 U1024 ( .B(n7395), .A(n4140), .S(n4152), .Y(n4986) );
  INVX1 U1025 ( .A(N4060), .Y(n7395) );
  MUX2X1 U1026 ( .B(n7394), .A(n4132), .S(n4152), .Y(n4985) );
  INVX1 U1027 ( .A(N4081), .Y(n7394) );
  MUX2X1 U1028 ( .B(n7346), .A(n4132), .S(n4153), .Y(n4984) );
  INVX1 U1029 ( .A(N4057), .Y(n7346) );
  MUX2X1 U1030 ( .B(n7347), .A(n4134), .S(n4153), .Y(n4983) );
  INVX1 U1031 ( .A(N4054), .Y(n7347) );
  MUX2X1 U1032 ( .B(n7348), .A(n4135), .S(n4153), .Y(n4982) );
  INVX1 U1033 ( .A(N4051), .Y(n7348) );
  MUX2X1 U1034 ( .B(n7349), .A(n4136), .S(n4153), .Y(n4981) );
  INVX1 U1035 ( .A(N4048), .Y(n7349) );
  MUX2X1 U1036 ( .B(n7350), .A(n4137), .S(n4153), .Y(n4980) );
  INVX1 U1037 ( .A(N4045), .Y(n7350) );
  MUX2X1 U1038 ( .B(n7351), .A(n4138), .S(n4153), .Y(n4979) );
  INVX1 U1039 ( .A(N4042), .Y(n7351) );
  MUX2X1 U1040 ( .B(n7352), .A(n4139), .S(n4153), .Y(n4978) );
  INVX1 U1041 ( .A(N4039), .Y(n7352) );
  MUX2X1 U1042 ( .B(n7353), .A(n4140), .S(n4153), .Y(n4977) );
  INVX1 U1043 ( .A(N4036), .Y(n7353) );
  MUX2X1 U1044 ( .B(n7330), .A(n4132), .S(n4154), .Y(n4976) );
  INVX1 U1045 ( .A(N4033), .Y(n7330) );
  MUX2X1 U1046 ( .B(n7331), .A(n4134), .S(n4154), .Y(n4975) );
  INVX1 U1047 ( .A(N4030), .Y(n7331) );
  MUX2X1 U1048 ( .B(n7332), .A(n4135), .S(n4154), .Y(n4974) );
  INVX1 U1049 ( .A(N4027), .Y(n7332) );
  MUX2X1 U1050 ( .B(n7333), .A(n4136), .S(n4154), .Y(n4973) );
  INVX1 U1051 ( .A(N4024), .Y(n7333) );
  MUX2X1 U1052 ( .B(n7334), .A(n4137), .S(n4154), .Y(n4972) );
  INVX1 U1053 ( .A(N4021), .Y(n7334) );
  MUX2X1 U1054 ( .B(n7335), .A(n4138), .S(n4154), .Y(n4971) );
  INVX1 U1055 ( .A(N4018), .Y(n7335) );
  MUX2X1 U1056 ( .B(n7336), .A(n4139), .S(n4154), .Y(n4970) );
  INVX1 U1057 ( .A(N4015), .Y(n7336) );
  MUX2X1 U1058 ( .B(n7337), .A(n4140), .S(n4154), .Y(n4969) );
  INVX1 U1059 ( .A(N4012), .Y(n7337) );
  MUX2X1 U1060 ( .B(n7577), .A(n4132), .S(n4155), .Y(n4968) );
  INVX1 U1061 ( .A(N4009), .Y(n7577) );
  MUX2X1 U1062 ( .B(n7576), .A(n4134), .S(n4155), .Y(n4967) );
  INVX1 U1063 ( .A(N4006), .Y(n7576) );
  MUX2X1 U1064 ( .B(n7575), .A(n4135), .S(n4155), .Y(n4966) );
  INVX1 U1065 ( .A(N4003), .Y(n7575) );
  MUX2X1 U1066 ( .B(n7574), .A(n4136), .S(n4155), .Y(n4965) );
  INVX1 U1067 ( .A(N4000), .Y(n7574) );
  MUX2X1 U1068 ( .B(n7573), .A(n4137), .S(n4155), .Y(n4964) );
  INVX1 U1069 ( .A(N3997), .Y(n7573) );
  MUX2X1 U1070 ( .B(n7572), .A(n4138), .S(n4155), .Y(n4963) );
  INVX1 U1071 ( .A(N3994), .Y(n7572) );
  MUX2X1 U1072 ( .B(n7571), .A(n4139), .S(n4155), .Y(n4962) );
  INVX1 U1073 ( .A(N3991), .Y(n7571) );
  MUX2X1 U1074 ( .B(n7570), .A(n4140), .S(n4155), .Y(n4961) );
  INVX1 U1075 ( .A(N3988), .Y(n7570) );
  MUX2X1 U1076 ( .B(n7593), .A(n4132), .S(n4156), .Y(n4960) );
  INVX1 U1077 ( .A(N3985), .Y(n7593) );
  MUX2X1 U1078 ( .B(n7592), .A(n4134), .S(n4156), .Y(n4959) );
  INVX1 U1079 ( .A(N3982), .Y(n7592) );
  MUX2X1 U1080 ( .B(n7591), .A(n4135), .S(n4156), .Y(n4958) );
  INVX1 U1081 ( .A(N3979), .Y(n7591) );
  MUX2X1 U1082 ( .B(n7590), .A(n4136), .S(n4156), .Y(n4957) );
  INVX1 U1083 ( .A(N3976), .Y(n7590) );
  MUX2X1 U1084 ( .B(n7589), .A(n4137), .S(n4156), .Y(n4956) );
  INVX1 U1085 ( .A(N3973), .Y(n7589) );
  MUX2X1 U1086 ( .B(n7588), .A(n4138), .S(n4156), .Y(n4955) );
  INVX1 U1087 ( .A(N3970), .Y(n7588) );
  MUX2X1 U1088 ( .B(n7587), .A(n4139), .S(n4156), .Y(n4954) );
  INVX1 U1089 ( .A(N3967), .Y(n7587) );
  MUX2X1 U1090 ( .B(n7586), .A(n4140), .S(n4156), .Y(n4953) );
  INVX1 U1091 ( .A(N3964), .Y(n7586) );
  MUX2X1 U1092 ( .B(n7609), .A(n4132), .S(n4157), .Y(n4952) );
  INVX1 U1093 ( .A(N3961), .Y(n7609) );
  MUX2X1 U1094 ( .B(n7608), .A(n4134), .S(n4157), .Y(n4951) );
  INVX1 U1095 ( .A(N3958), .Y(n7608) );
  MUX2X1 U1096 ( .B(n7607), .A(n4135), .S(n4157), .Y(n4950) );
  INVX1 U1097 ( .A(N3955), .Y(n7607) );
  MUX2X1 U1098 ( .B(n7606), .A(n4136), .S(n4157), .Y(n4949) );
  INVX1 U1099 ( .A(N3952), .Y(n7606) );
  MUX2X1 U1100 ( .B(n7605), .A(n4137), .S(n4157), .Y(n4948) );
  INVX1 U1101 ( .A(N3949), .Y(n7605) );
  MUX2X1 U1102 ( .B(n7604), .A(n4138), .S(n4157), .Y(n4947) );
  INVX1 U1103 ( .A(N3946), .Y(n7604) );
  MUX2X1 U1104 ( .B(n7603), .A(n4139), .S(n4157), .Y(n4946) );
  INVX1 U1105 ( .A(N3943), .Y(n7603) );
  MUX2X1 U1106 ( .B(n7602), .A(n4140), .S(n4157), .Y(n4945) );
  INVX1 U1107 ( .A(N3940), .Y(n7602) );
  MUX2X1 U1108 ( .B(n7625), .A(n4132), .S(n4158), .Y(n4944) );
  INVX1 U1109 ( .A(N3937), .Y(n7625) );
  MUX2X1 U1110 ( .B(n7624), .A(n4134), .S(n4158), .Y(n4943) );
  INVX1 U1111 ( .A(N3934), .Y(n7624) );
  MUX2X1 U1112 ( .B(n7623), .A(n4135), .S(n4158), .Y(n4942) );
  INVX1 U1113 ( .A(N3931), .Y(n7623) );
  MUX2X1 U1114 ( .B(n7622), .A(n4136), .S(n4158), .Y(n4941) );
  INVX1 U1115 ( .A(N3928), .Y(n7622) );
  MUX2X1 U1116 ( .B(n7621), .A(n4137), .S(n4158), .Y(n4940) );
  INVX1 U1117 ( .A(N3925), .Y(n7621) );
  MUX2X1 U1118 ( .B(n7620), .A(n4138), .S(n4158), .Y(n4939) );
  INVX1 U1119 ( .A(N3922), .Y(n7620) );
  MUX2X1 U1120 ( .B(n7619), .A(n4139), .S(n4158), .Y(n4938) );
  INVX1 U1121 ( .A(N3919), .Y(n7619) );
  MUX2X1 U1122 ( .B(n7618), .A(n4140), .S(n4158), .Y(n4937) );
  INVX1 U1123 ( .A(N3916), .Y(n7618) );
  MUX2X1 U1124 ( .B(n7641), .A(n4132), .S(n4159), .Y(n4936) );
  INVX1 U1125 ( .A(N3913), .Y(n7641) );
  MUX2X1 U1126 ( .B(n7640), .A(n4134), .S(n4159), .Y(n4935) );
  INVX1 U1127 ( .A(N3910), .Y(n7640) );
  MUX2X1 U1128 ( .B(n7639), .A(n4135), .S(n4159), .Y(n4934) );
  INVX1 U1129 ( .A(N3907), .Y(n7639) );
  MUX2X1 U1130 ( .B(n7638), .A(n4136), .S(n4159), .Y(n4933) );
  INVX1 U1131 ( .A(N3904), .Y(n7638) );
  MUX2X1 U1132 ( .B(n7637), .A(n4137), .S(n4159), .Y(n4932) );
  INVX1 U1133 ( .A(N3901), .Y(n7637) );
  MUX2X1 U1134 ( .B(n7636), .A(n4138), .S(n4159), .Y(n4931) );
  INVX1 U1135 ( .A(N3898), .Y(n7636) );
  MUX2X1 U1136 ( .B(n7635), .A(n4139), .S(n4159), .Y(n4930) );
  INVX1 U1137 ( .A(N3895), .Y(n7635) );
  MUX2X1 U1138 ( .B(n7634), .A(n4140), .S(n4159), .Y(n4929) );
  INVX1 U1139 ( .A(N3892), .Y(n7634) );
  MUX2X1 U1140 ( .B(n7657), .A(n4132), .S(n4160), .Y(n4928) );
  INVX1 U1141 ( .A(N3889), .Y(n7657) );
  MUX2X1 U1142 ( .B(n7656), .A(n4134), .S(n4160), .Y(n4927) );
  INVX1 U1143 ( .A(N3886), .Y(n7656) );
  MUX2X1 U1144 ( .B(n7655), .A(n4135), .S(n4160), .Y(n4926) );
  INVX1 U1145 ( .A(N3883), .Y(n7655) );
  MUX2X1 U1146 ( .B(n7654), .A(n4136), .S(n4160), .Y(n4925) );
  INVX1 U1147 ( .A(N3880), .Y(n7654) );
  MUX2X1 U1148 ( .B(n7653), .A(n4137), .S(n4160), .Y(n4924) );
  INVX1 U1149 ( .A(N3877), .Y(n7653) );
  MUX2X1 U1150 ( .B(n7652), .A(n4138), .S(n4160), .Y(n4923) );
  INVX1 U1151 ( .A(N3874), .Y(n7652) );
  MUX2X1 U1152 ( .B(n7651), .A(n4139), .S(n4160), .Y(n4922) );
  INVX1 U1153 ( .A(N3871), .Y(n7651) );
  MUX2X1 U1154 ( .B(n7650), .A(n4140), .S(n4160), .Y(n4921) );
  INVX1 U1155 ( .A(N3868), .Y(n7650) );
  MUX2X1 U1156 ( .B(n7673), .A(n4132), .S(n4161), .Y(n4920) );
  INVX1 U1157 ( .A(N3865), .Y(n7673) );
  MUX2X1 U1158 ( .B(n7672), .A(n4134), .S(n4161), .Y(n4919) );
  INVX1 U1159 ( .A(N3862), .Y(n7672) );
  MUX2X1 U1160 ( .B(n7671), .A(n4135), .S(n4161), .Y(n4918) );
  INVX1 U1161 ( .A(N3859), .Y(n7671) );
  MUX2X1 U1162 ( .B(n7670), .A(n4136), .S(n4161), .Y(n4917) );
  INVX1 U1163 ( .A(N3856), .Y(n7670) );
  MUX2X1 U1164 ( .B(n7669), .A(n4137), .S(n4161), .Y(n4916) );
  INVX1 U1165 ( .A(N3853), .Y(n7669) );
  MUX2X1 U1166 ( .B(n7668), .A(n4138), .S(n4161), .Y(n4915) );
  INVX1 U1167 ( .A(N3850), .Y(n7668) );
  MUX2X1 U1168 ( .B(n7667), .A(n4139), .S(n4161), .Y(n4914) );
  INVX1 U1169 ( .A(N3847), .Y(n7667) );
  MUX2X1 U1170 ( .B(n7666), .A(n4140), .S(n4161), .Y(n4913) );
  INVX1 U1171 ( .A(N3844), .Y(n7666) );
  MUX2X1 U1172 ( .B(n7321), .A(n4132), .S(n4162), .Y(n4912) );
  INVX1 U1173 ( .A(N3841), .Y(n7321) );
  MUX2X1 U1174 ( .B(n7320), .A(n4134), .S(n4162), .Y(n4911) );
  INVX1 U1175 ( .A(N3838), .Y(n7320) );
  MUX2X1 U1176 ( .B(n7319), .A(n4135), .S(n4162), .Y(n4910) );
  INVX1 U1177 ( .A(N3835), .Y(n7319) );
  MUX2X1 U1178 ( .B(n7318), .A(n4136), .S(n4162), .Y(n4909) );
  INVX1 U1179 ( .A(N3832), .Y(n7318) );
  MUX2X1 U1180 ( .B(n7317), .A(n4137), .S(n4162), .Y(n4908) );
  INVX1 U1181 ( .A(N3829), .Y(n7317) );
  MUX2X1 U1182 ( .B(n7316), .A(n4138), .S(n4162), .Y(n4907) );
  INVX1 U1183 ( .A(N3826), .Y(n7316) );
  MUX2X1 U1184 ( .B(n7315), .A(n4139), .S(n4162), .Y(n4906) );
  INVX1 U1185 ( .A(N3823), .Y(n7315) );
  MUX2X1 U1186 ( .B(n7314), .A(n4140), .S(n4162), .Y(n4905) );
  INVX1 U1187 ( .A(N3820), .Y(n7314) );
  MUX2X1 U1188 ( .B(n7305), .A(n4132), .S(n4163), .Y(n4904) );
  INVX1 U1189 ( .A(N3817), .Y(n7305) );
  MUX2X1 U1190 ( .B(n7304), .A(n4134), .S(n4163), .Y(n4903) );
  INVX1 U1191 ( .A(N3814), .Y(n7304) );
  MUX2X1 U1192 ( .B(n7303), .A(n4135), .S(n4163), .Y(n4902) );
  INVX1 U1193 ( .A(N3811), .Y(n7303) );
  MUX2X1 U1194 ( .B(n7302), .A(n4136), .S(n4163), .Y(n4901) );
  INVX1 U1195 ( .A(N3808), .Y(n7302) );
  MUX2X1 U1196 ( .B(n7301), .A(n4137), .S(n4163), .Y(n4900) );
  INVX1 U1197 ( .A(N3805), .Y(n7301) );
  MUX2X1 U1198 ( .B(n7300), .A(n4138), .S(n4163), .Y(n4899) );
  INVX1 U1199 ( .A(N3802), .Y(n7300) );
  MUX2X1 U1200 ( .B(n7299), .A(n4139), .S(n4163), .Y(n4898) );
  INVX1 U1201 ( .A(N3799), .Y(n7299) );
  MUX2X1 U1202 ( .B(n7298), .A(n4140), .S(n4163), .Y(n4897) );
  INVX1 U1203 ( .A(N3796), .Y(n7298) );
  MUX2X1 U1204 ( .B(n7689), .A(n4137), .S(n4164), .Y(n4896) );
  NAND2X1 U1205 ( .A(n4165), .B(InData[4]), .Y(n4137) );
  INVX1 U1206 ( .A(N3781), .Y(n7689) );
  MUX2X1 U1207 ( .B(n7688), .A(n4138), .S(n4164), .Y(n4895) );
  NAND2X1 U1208 ( .A(n4165), .B(InData[5]), .Y(n4138) );
  INVX1 U1209 ( .A(N3778), .Y(n7688) );
  MUX2X1 U1210 ( .B(n7687), .A(n4139), .S(n4164), .Y(n4894) );
  NAND2X1 U1211 ( .A(n4165), .B(InData[6]), .Y(n4139) );
  INVX1 U1212 ( .A(N3775), .Y(n7687) );
  MUX2X1 U1213 ( .B(n7686), .A(n4140), .S(n4164), .Y(n4893) );
  NAND2X1 U1214 ( .A(n4165), .B(InData[7]), .Y(n4140) );
  INVX1 U1215 ( .A(N3772), .Y(n7686) );
  MUX2X1 U1216 ( .B(n7685), .A(n4132), .S(n4164), .Y(n4892) );
  NAND2X1 U1217 ( .A(n4165), .B(InData[0]), .Y(n4132) );
  INVX1 U1218 ( .A(N3793), .Y(n7685) );
  MUX2X1 U1219 ( .B(n7684), .A(n4134), .S(n4164), .Y(n4891) );
  NAND2X1 U1220 ( .A(n4165), .B(InData[1]), .Y(n4134) );
  INVX1 U1221 ( .A(N3790), .Y(n7684) );
  MUX2X1 U1222 ( .B(n7683), .A(n4135), .S(n4164), .Y(n4890) );
  NAND2X1 U1223 ( .A(n4165), .B(InData[2]), .Y(n4135) );
  INVX1 U1224 ( .A(N3787), .Y(n7683) );
  MUX2X1 U1225 ( .B(n7682), .A(n4136), .S(n4164), .Y(n4889) );
  NAND2X1 U1226 ( .A(n4165), .B(InData[3]), .Y(n4136) );
  INVX1 U1227 ( .A(n4166), .Y(n4165) );
  INVX1 U1228 ( .A(N3784), .Y(n7682) );
  OAI21X1 U1229 ( .A(n7530), .B(n4133), .C(n4167), .Y(n4888) );
  INVX1 U1230 ( .A(N4370), .Y(n7530) );
  OAI21X1 U1231 ( .A(n7531), .B(n4133), .C(n4167), .Y(n4887) );
  INVX1 U1232 ( .A(N4367), .Y(n7531) );
  OAI21X1 U1233 ( .A(n7532), .B(n4133), .C(n4167), .Y(n4886) );
  INVX1 U1234 ( .A(N4364), .Y(n7532) );
  OAI21X1 U1235 ( .A(n7533), .B(n4133), .C(n4167), .Y(n4885) );
  INVX1 U1236 ( .A(N4361), .Y(n7533) );
  OAI21X1 U1237 ( .A(n7534), .B(n4133), .C(n4167), .Y(n4884) );
  INVX1 U1238 ( .A(N4358), .Y(n7534) );
  OAI21X1 U1239 ( .A(n7535), .B(n4133), .C(n4167), .Y(n4883) );
  INVX1 U1240 ( .A(N4355), .Y(n7535) );
  OAI21X1 U1241 ( .A(n7536), .B(n4133), .C(n4167), .Y(n4882) );
  INVX1 U1242 ( .A(N4352), .Y(n7536) );
  OAI21X1 U1243 ( .A(n7537), .B(n4133), .C(n4167), .Y(n4881) );
  NAND2X1 U1244 ( .A(n4168), .B(n4133), .Y(n4167) );
  INVX1 U1245 ( .A(n4169), .Y(n4133) );
  NAND3X1 U1246 ( .A(n3582), .B(n3580), .C(n4170), .Y(n4169) );
  INVX1 U1247 ( .A(N4349), .Y(n7537) );
  OAI21X1 U1248 ( .A(n7521), .B(n4141), .C(n4171), .Y(n4880) );
  INVX1 U1249 ( .A(N4346), .Y(n7521) );
  OAI21X1 U1250 ( .A(n7520), .B(n4141), .C(n4171), .Y(n4879) );
  INVX1 U1251 ( .A(N4343), .Y(n7520) );
  OAI21X1 U1252 ( .A(n7519), .B(n4141), .C(n4171), .Y(n4878) );
  INVX1 U1253 ( .A(N4340), .Y(n7519) );
  OAI21X1 U1254 ( .A(n7518), .B(n4141), .C(n4171), .Y(n4877) );
  INVX1 U1255 ( .A(N4337), .Y(n7518) );
  OAI21X1 U1256 ( .A(n7517), .B(n4141), .C(n4171), .Y(n4876) );
  INVX1 U1257 ( .A(N4334), .Y(n7517) );
  OAI21X1 U1258 ( .A(n7516), .B(n4141), .C(n4171), .Y(n4875) );
  INVX1 U1259 ( .A(N4331), .Y(n7516) );
  OAI21X1 U1260 ( .A(n7515), .B(n4141), .C(n4171), .Y(n4874) );
  INVX1 U1261 ( .A(N4328), .Y(n7515) );
  OAI21X1 U1262 ( .A(n7514), .B(n4141), .C(n4171), .Y(n4873) );
  NAND2X1 U1263 ( .A(n4168), .B(n4141), .Y(n4171) );
  AND2X1 U1264 ( .A(n4172), .B(n4173), .Y(n4141) );
  INVX1 U1265 ( .A(N4325), .Y(n7514) );
  OAI21X1 U1266 ( .A(n7505), .B(n4142), .C(n4174), .Y(n4872) );
  INVX1 U1267 ( .A(N4322), .Y(n7505) );
  OAI21X1 U1268 ( .A(n7504), .B(n4142), .C(n4174), .Y(n4871) );
  INVX1 U1269 ( .A(N4319), .Y(n7504) );
  OAI21X1 U1270 ( .A(n7503), .B(n4142), .C(n4174), .Y(n4870) );
  INVX1 U1271 ( .A(N4316), .Y(n7503) );
  OAI21X1 U1272 ( .A(n7502), .B(n4142), .C(n4174), .Y(n4869) );
  INVX1 U1273 ( .A(N4313), .Y(n7502) );
  OAI21X1 U1274 ( .A(n7501), .B(n4142), .C(n4174), .Y(n4868) );
  INVX1 U1275 ( .A(N4310), .Y(n7501) );
  OAI21X1 U1276 ( .A(n7500), .B(n4142), .C(n4174), .Y(n4867) );
  INVX1 U1277 ( .A(N4307), .Y(n7500) );
  OAI21X1 U1278 ( .A(n7499), .B(n4142), .C(n4174), .Y(n4866) );
  INVX1 U1279 ( .A(N4304), .Y(n7499) );
  OAI21X1 U1280 ( .A(n7498), .B(n4142), .C(n4174), .Y(n4865) );
  NAND2X1 U1281 ( .A(n4168), .B(n4142), .Y(n4174) );
  AND2X1 U1282 ( .A(n4172), .B(n4175), .Y(n4142) );
  INVX1 U1283 ( .A(N4301), .Y(n7498) );
  OAI21X1 U1284 ( .A(n7457), .B(n4143), .C(n4176), .Y(n4864) );
  INVX1 U1285 ( .A(N4298), .Y(n7457) );
  OAI21X1 U1286 ( .A(n7456), .B(n4143), .C(n4176), .Y(n4863) );
  INVX1 U1287 ( .A(N4295), .Y(n7456) );
  OAI21X1 U1288 ( .A(n7455), .B(n4143), .C(n4176), .Y(n4862) );
  INVX1 U1289 ( .A(N4292), .Y(n7455) );
  OAI21X1 U1290 ( .A(n7454), .B(n4143), .C(n4176), .Y(n4861) );
  INVX1 U1291 ( .A(N4289), .Y(n7454) );
  OAI21X1 U1292 ( .A(n7453), .B(n4143), .C(n4176), .Y(n4860) );
  INVX1 U1293 ( .A(N4286), .Y(n7453) );
  OAI21X1 U1294 ( .A(n7452), .B(n4143), .C(n4176), .Y(n4859) );
  INVX1 U1295 ( .A(N4283), .Y(n7452) );
  OAI21X1 U1296 ( .A(n7451), .B(n4143), .C(n4176), .Y(n4858) );
  INVX1 U1297 ( .A(N4280), .Y(n7451) );
  OAI21X1 U1298 ( .A(n7450), .B(n4143), .C(n4176), .Y(n4857) );
  NAND2X1 U1299 ( .A(n4168), .B(n4143), .Y(n4176) );
  AND2X1 U1300 ( .A(n4177), .B(n4173), .Y(n4143) );
  INVX1 U1301 ( .A(N4277), .Y(n7450) );
  OAI21X1 U1302 ( .A(n7441), .B(n4144), .C(n4178), .Y(n4856) );
  INVX1 U1303 ( .A(N4274), .Y(n7441) );
  OAI21X1 U1304 ( .A(n7440), .B(n4144), .C(n4178), .Y(n4855) );
  INVX1 U1305 ( .A(N4271), .Y(n7440) );
  OAI21X1 U1306 ( .A(n7439), .B(n4144), .C(n4178), .Y(n4854) );
  INVX1 U1307 ( .A(N4268), .Y(n7439) );
  OAI21X1 U1308 ( .A(n7438), .B(n4144), .C(n4178), .Y(n4853) );
  INVX1 U1309 ( .A(N4265), .Y(n7438) );
  OAI21X1 U1310 ( .A(n7437), .B(n4144), .C(n4178), .Y(n4852) );
  INVX1 U1311 ( .A(N4262), .Y(n7437) );
  OAI21X1 U1312 ( .A(n7436), .B(n4144), .C(n4178), .Y(n4851) );
  INVX1 U1313 ( .A(N4259), .Y(n7436) );
  OAI21X1 U1314 ( .A(n7435), .B(n4144), .C(n4178), .Y(n4850) );
  INVX1 U1315 ( .A(N4256), .Y(n7435) );
  OAI21X1 U1316 ( .A(n7434), .B(n4144), .C(n4178), .Y(n4849) );
  NAND2X1 U1317 ( .A(n4168), .B(n4144), .Y(n4178) );
  AND2X1 U1318 ( .A(n4177), .B(n4175), .Y(n4144) );
  INVX1 U1319 ( .A(N4253), .Y(n7434) );
  OAI21X1 U1320 ( .A(n7393), .B(n4145), .C(n4179), .Y(n4848) );
  INVX1 U1321 ( .A(N4250), .Y(n7393) );
  OAI21X1 U1322 ( .A(n7392), .B(n4145), .C(n4179), .Y(n4847) );
  INVX1 U1323 ( .A(N4247), .Y(n7392) );
  OAI21X1 U1324 ( .A(n7391), .B(n4145), .C(n4179), .Y(n4846) );
  INVX1 U1325 ( .A(N4244), .Y(n7391) );
  OAI21X1 U1326 ( .A(n7390), .B(n4145), .C(n4179), .Y(n4845) );
  INVX1 U1327 ( .A(N4241), .Y(n7390) );
  OAI21X1 U1328 ( .A(n7389), .B(n4145), .C(n4179), .Y(n4844) );
  INVX1 U1329 ( .A(N4238), .Y(n7389) );
  OAI21X1 U1330 ( .A(n7388), .B(n4145), .C(n4179), .Y(n4843) );
  INVX1 U1331 ( .A(N4235), .Y(n7388) );
  OAI21X1 U1332 ( .A(n7387), .B(n4145), .C(n4179), .Y(n4842) );
  INVX1 U1333 ( .A(N4232), .Y(n7387) );
  OAI21X1 U1334 ( .A(n7386), .B(n4145), .C(n4179), .Y(n4841) );
  NAND2X1 U1335 ( .A(n4168), .B(n4145), .Y(n4179) );
  AND2X1 U1336 ( .A(n4180), .B(n4173), .Y(n4145) );
  INVX1 U1337 ( .A(n3598), .Y(n4173) );
  NAND2X1 U1338 ( .A(n4181), .B(n3664), .Y(n3598) );
  INVX1 U1339 ( .A(N4229), .Y(n7386) );
  OAI21X1 U1340 ( .A(n7377), .B(n4146), .C(n4182), .Y(n4840) );
  INVX1 U1341 ( .A(N4226), .Y(n7377) );
  OAI21X1 U1342 ( .A(n7376), .B(n4146), .C(n4182), .Y(n4839) );
  INVX1 U1343 ( .A(N4223), .Y(n7376) );
  OAI21X1 U1344 ( .A(n7375), .B(n4146), .C(n4182), .Y(n4838) );
  INVX1 U1345 ( .A(N4220), .Y(n7375) );
  OAI21X1 U1346 ( .A(n7374), .B(n4146), .C(n4182), .Y(n4837) );
  INVX1 U1347 ( .A(N4217), .Y(n7374) );
  OAI21X1 U1348 ( .A(n7373), .B(n4146), .C(n4182), .Y(n4836) );
  INVX1 U1349 ( .A(N4214), .Y(n7373) );
  OAI21X1 U1350 ( .A(n7372), .B(n4146), .C(n4182), .Y(n4835) );
  INVX1 U1351 ( .A(N4211), .Y(n7372) );
  OAI21X1 U1352 ( .A(n7371), .B(n4146), .C(n4182), .Y(n4834) );
  INVX1 U1353 ( .A(N4208), .Y(n7371) );
  OAI21X1 U1354 ( .A(n7370), .B(n4146), .C(n4182), .Y(n4833) );
  NAND2X1 U1355 ( .A(n4168), .B(n4146), .Y(n4182) );
  AND2X1 U1356 ( .A(n4180), .B(n4175), .Y(n4146) );
  INVX1 U1357 ( .A(n3610), .Y(n4175) );
  NAND2X1 U1358 ( .A(n4183), .B(n3664), .Y(n3610) );
  INVX1 U1359 ( .A(N4205), .Y(n7370) );
  OAI21X1 U1360 ( .A(n7546), .B(n4147), .C(n4184), .Y(n4832) );
  INVX1 U1361 ( .A(N4202), .Y(n7546) );
  OAI21X1 U1362 ( .A(n7547), .B(n4147), .C(n4184), .Y(n4831) );
  INVX1 U1363 ( .A(N4199), .Y(n7547) );
  OAI21X1 U1364 ( .A(n7548), .B(n4147), .C(n4184), .Y(n4830) );
  INVX1 U1365 ( .A(N4196), .Y(n7548) );
  OAI21X1 U1366 ( .A(n7549), .B(n4147), .C(n4184), .Y(n4829) );
  INVX1 U1367 ( .A(N4193), .Y(n7549) );
  OAI21X1 U1368 ( .A(n7550), .B(n4147), .C(n4184), .Y(n4828) );
  INVX1 U1369 ( .A(N4190), .Y(n7550) );
  OAI21X1 U1370 ( .A(n7551), .B(n4147), .C(n4184), .Y(n4827) );
  INVX1 U1371 ( .A(N4187), .Y(n7551) );
  OAI21X1 U1372 ( .A(n7552), .B(n4147), .C(n4184), .Y(n4826) );
  INVX1 U1373 ( .A(N4184), .Y(n7552) );
  OAI21X1 U1374 ( .A(n7553), .B(n4147), .C(n4184), .Y(n4825) );
  NAND2X1 U1375 ( .A(n4168), .B(n4147), .Y(n4184) );
  INVX1 U1376 ( .A(n4185), .Y(n4147) );
  NAND3X1 U1377 ( .A(n3665), .B(n3664), .C(n4170), .Y(n4185) );
  INVX1 U1378 ( .A(N4181), .Y(n7553) );
  OAI21X1 U1379 ( .A(n7562), .B(n4148), .C(n4186), .Y(n4824) );
  INVX1 U1380 ( .A(N4178), .Y(n7562) );
  OAI21X1 U1381 ( .A(n7563), .B(n4148), .C(n4186), .Y(n4823) );
  INVX1 U1382 ( .A(N4175), .Y(n7563) );
  OAI21X1 U1383 ( .A(n7564), .B(n4148), .C(n4186), .Y(n4822) );
  INVX1 U1384 ( .A(N4172), .Y(n7564) );
  OAI21X1 U1385 ( .A(n7565), .B(n4148), .C(n4186), .Y(n4821) );
  INVX1 U1386 ( .A(N4169), .Y(n7565) );
  OAI21X1 U1387 ( .A(n7566), .B(n4148), .C(n4186), .Y(n4820) );
  INVX1 U1388 ( .A(N4166), .Y(n7566) );
  OAI21X1 U1389 ( .A(n7567), .B(n4148), .C(n4186), .Y(n4819) );
  INVX1 U1390 ( .A(N4163), .Y(n7567) );
  OAI21X1 U1391 ( .A(n7568), .B(n4148), .C(n4186), .Y(n4818) );
  INVX1 U1392 ( .A(N4160), .Y(n7568) );
  OAI21X1 U1393 ( .A(n7569), .B(n4148), .C(n4186), .Y(n4817) );
  NAND2X1 U1394 ( .A(n4168), .B(n4148), .Y(n4186) );
  NOR2X1 U1395 ( .A(n4187), .B(n3676), .Y(n4148) );
  INVX1 U1396 ( .A(N4157), .Y(n7569) );
  OAI21X1 U1397 ( .A(n7489), .B(n4149), .C(n4188), .Y(n4816) );
  INVX1 U1398 ( .A(N4154), .Y(n7489) );
  OAI21X1 U1399 ( .A(n7488), .B(n4149), .C(n4188), .Y(n4815) );
  INVX1 U1400 ( .A(N4151), .Y(n7488) );
  OAI21X1 U1401 ( .A(n7487), .B(n4149), .C(n4188), .Y(n4814) );
  INVX1 U1402 ( .A(N4148), .Y(n7487) );
  OAI21X1 U1403 ( .A(n7486), .B(n4149), .C(n4188), .Y(n4813) );
  INVX1 U1404 ( .A(N4145), .Y(n7486) );
  OAI21X1 U1405 ( .A(n7485), .B(n4149), .C(n4188), .Y(n4812) );
  INVX1 U1406 ( .A(N4142), .Y(n7485) );
  OAI21X1 U1407 ( .A(n7484), .B(n4149), .C(n4188), .Y(n4811) );
  INVX1 U1408 ( .A(N4139), .Y(n7484) );
  OAI21X1 U1409 ( .A(n7483), .B(n4149), .C(n4188), .Y(n4810) );
  INVX1 U1410 ( .A(N4136), .Y(n7483) );
  OAI21X1 U1411 ( .A(n7482), .B(n4149), .C(n4188), .Y(n4809) );
  NAND2X1 U1412 ( .A(n4168), .B(n4149), .Y(n4188) );
  AND2X1 U1413 ( .A(n4172), .B(n4189), .Y(n4149) );
  INVX1 U1414 ( .A(N4133), .Y(n7482) );
  OAI21X1 U1415 ( .A(n7473), .B(n4150), .C(n4190), .Y(n4808) );
  INVX1 U1416 ( .A(N4130), .Y(n7473) );
  OAI21X1 U1417 ( .A(n7472), .B(n4150), .C(n4190), .Y(n4807) );
  INVX1 U1418 ( .A(N4127), .Y(n7472) );
  OAI21X1 U1419 ( .A(n7471), .B(n4150), .C(n4190), .Y(n4806) );
  INVX1 U1420 ( .A(N4124), .Y(n7471) );
  OAI21X1 U1421 ( .A(n7470), .B(n4150), .C(n4190), .Y(n4805) );
  INVX1 U1422 ( .A(N4121), .Y(n7470) );
  OAI21X1 U1423 ( .A(n7469), .B(n4150), .C(n4190), .Y(n4804) );
  INVX1 U1424 ( .A(N4118), .Y(n7469) );
  OAI21X1 U1425 ( .A(n7468), .B(n4150), .C(n4190), .Y(n4803) );
  INVX1 U1426 ( .A(N4115), .Y(n7468) );
  OAI21X1 U1427 ( .A(n7467), .B(n4150), .C(n4190), .Y(n4802) );
  INVX1 U1428 ( .A(N4112), .Y(n7467) );
  OAI21X1 U1429 ( .A(n7466), .B(n4150), .C(n4190), .Y(n4801) );
  NAND2X1 U1430 ( .A(n4168), .B(n4150), .Y(n4190) );
  AND2X1 U1431 ( .A(n4172), .B(n4191), .Y(n4150) );
  AND2X1 U1432 ( .A(n4170), .B(n3766), .Y(n4172) );
  INVX1 U1433 ( .A(N4109), .Y(n7466) );
  OAI21X1 U1434 ( .A(n7425), .B(n4151), .C(n4192), .Y(n4800) );
  INVX1 U1435 ( .A(N4106), .Y(n7425) );
  OAI21X1 U1436 ( .A(n7424), .B(n4151), .C(n4192), .Y(n4799) );
  INVX1 U1437 ( .A(N4103), .Y(n7424) );
  OAI21X1 U1438 ( .A(n7423), .B(n4151), .C(n4192), .Y(n4798) );
  INVX1 U1439 ( .A(N4100), .Y(n7423) );
  OAI21X1 U1440 ( .A(n7422), .B(n4151), .C(n4192), .Y(n4797) );
  INVX1 U1441 ( .A(N4097), .Y(n7422) );
  OAI21X1 U1442 ( .A(n7421), .B(n4151), .C(n4192), .Y(n4796) );
  INVX1 U1443 ( .A(N4094), .Y(n7421) );
  OAI21X1 U1444 ( .A(n7420), .B(n4151), .C(n4192), .Y(n4795) );
  INVX1 U1445 ( .A(N4091), .Y(n7420) );
  OAI21X1 U1446 ( .A(n7419), .B(n4151), .C(n4192), .Y(n4794) );
  INVX1 U1447 ( .A(N4088), .Y(n7419) );
  OAI21X1 U1448 ( .A(n7418), .B(n4151), .C(n4192), .Y(n4793) );
  NAND2X1 U1449 ( .A(n4168), .B(n4151), .Y(n4192) );
  AND2X1 U1450 ( .A(n4177), .B(n4189), .Y(n4151) );
  INVX1 U1451 ( .A(N4085), .Y(n7418) );
  OAI21X1 U1452 ( .A(n7402), .B(n4152), .C(n4193), .Y(n4792) );
  INVX1 U1453 ( .A(N4082), .Y(n7402) );
  OAI21X1 U1454 ( .A(n7403), .B(n4152), .C(n4193), .Y(n4791) );
  INVX1 U1455 ( .A(N4079), .Y(n7403) );
  OAI21X1 U1456 ( .A(n7404), .B(n4152), .C(n4193), .Y(n4790) );
  INVX1 U1457 ( .A(N4076), .Y(n7404) );
  OAI21X1 U1458 ( .A(n7405), .B(n4152), .C(n4193), .Y(n4789) );
  INVX1 U1459 ( .A(N4073), .Y(n7405) );
  OAI21X1 U1460 ( .A(n7406), .B(n4152), .C(n4193), .Y(n4788) );
  INVX1 U1461 ( .A(N4070), .Y(n7406) );
  OAI21X1 U1462 ( .A(n7407), .B(n4152), .C(n4193), .Y(n4787) );
  INVX1 U1463 ( .A(N4067), .Y(n7407) );
  OAI21X1 U1464 ( .A(n7408), .B(n4152), .C(n4193), .Y(n4786) );
  INVX1 U1465 ( .A(N4064), .Y(n7408) );
  OAI21X1 U1466 ( .A(n7409), .B(n4152), .C(n4193), .Y(n4785) );
  NAND2X1 U1467 ( .A(n4168), .B(n4152), .Y(n4193) );
  AND2X1 U1468 ( .A(n4177), .B(n4191), .Y(n4152) );
  AND2X1 U1469 ( .A(n4170), .B(n3785), .Y(n4177) );
  INVX1 U1470 ( .A(N4061), .Y(n7409) );
  OAI21X1 U1471 ( .A(n7361), .B(n4153), .C(n4194), .Y(n4784) );
  INVX1 U1472 ( .A(N4058), .Y(n7361) );
  OAI21X1 U1473 ( .A(n7360), .B(n4153), .C(n4194), .Y(n4783) );
  INVX1 U1474 ( .A(N4055), .Y(n7360) );
  OAI21X1 U1475 ( .A(n7359), .B(n4153), .C(n4194), .Y(n4782) );
  INVX1 U1476 ( .A(N4052), .Y(n7359) );
  OAI21X1 U1477 ( .A(n7358), .B(n4153), .C(n4194), .Y(n4781) );
  INVX1 U1478 ( .A(N4049), .Y(n7358) );
  OAI21X1 U1479 ( .A(n7357), .B(n4153), .C(n4194), .Y(n4780) );
  INVX1 U1480 ( .A(N4046), .Y(n7357) );
  OAI21X1 U1481 ( .A(n7356), .B(n4153), .C(n4194), .Y(n4779) );
  INVX1 U1482 ( .A(N4043), .Y(n7356) );
  OAI21X1 U1483 ( .A(n7355), .B(n4153), .C(n4194), .Y(n4778) );
  INVX1 U1484 ( .A(N4040), .Y(n7355) );
  OAI21X1 U1485 ( .A(n7354), .B(n4153), .C(n4194), .Y(n4777) );
  NAND2X1 U1486 ( .A(n4168), .B(n4153), .Y(n4194) );
  AND2X1 U1487 ( .A(n4180), .B(n4189), .Y(n4153) );
  INVX1 U1488 ( .A(n3755), .Y(n4189) );
  NAND2X1 U1489 ( .A(n4195), .B(n3815), .Y(n3755) );
  INVX1 U1490 ( .A(N4037), .Y(n7354) );
  OAI21X1 U1491 ( .A(n7345), .B(n4154), .C(n4196), .Y(n4776) );
  INVX1 U1492 ( .A(N4034), .Y(n7345) );
  OAI21X1 U1493 ( .A(n7344), .B(n4154), .C(n4196), .Y(n4775) );
  INVX1 U1494 ( .A(N4031), .Y(n7344) );
  OAI21X1 U1495 ( .A(n7343), .B(n4154), .C(n4196), .Y(n4774) );
  INVX1 U1496 ( .A(N4028), .Y(n7343) );
  OAI21X1 U1497 ( .A(n7342), .B(n4154), .C(n4196), .Y(n4773) );
  INVX1 U1498 ( .A(N4025), .Y(n7342) );
  OAI21X1 U1499 ( .A(n7341), .B(n4154), .C(n4196), .Y(n4772) );
  INVX1 U1500 ( .A(N4022), .Y(n7341) );
  OAI21X1 U1501 ( .A(n7340), .B(n4154), .C(n4196), .Y(n4771) );
  INVX1 U1502 ( .A(N4019), .Y(n7340) );
  OAI21X1 U1503 ( .A(n7339), .B(n4154), .C(n4196), .Y(n4770) );
  INVX1 U1504 ( .A(N4016), .Y(n7339) );
  OAI21X1 U1505 ( .A(n7338), .B(n4154), .C(n4196), .Y(n4769) );
  NAND2X1 U1506 ( .A(n4168), .B(n4154), .Y(n4196) );
  AND2X1 U1507 ( .A(n4180), .B(n4191), .Y(n4154) );
  INVX1 U1508 ( .A(n3765), .Y(n4191) );
  NAND2X1 U1509 ( .A(n4197), .B(n3815), .Y(n3765) );
  AND2X1 U1510 ( .A(n4170), .B(n3804), .Y(n4180) );
  INVX1 U1511 ( .A(N4013), .Y(n7338) );
  OAI21X1 U1512 ( .A(n7578), .B(n4155), .C(n4198), .Y(n4768) );
  INVX1 U1513 ( .A(N4010), .Y(n7578) );
  OAI21X1 U1514 ( .A(n7579), .B(n4155), .C(n4198), .Y(n4767) );
  INVX1 U1515 ( .A(N4007), .Y(n7579) );
  OAI21X1 U1516 ( .A(n7580), .B(n4155), .C(n4198), .Y(n4766) );
  INVX1 U1517 ( .A(N4004), .Y(n7580) );
  OAI21X1 U1518 ( .A(n7581), .B(n4155), .C(n4198), .Y(n4765) );
  INVX1 U1519 ( .A(N4001), .Y(n7581) );
  OAI21X1 U1520 ( .A(n7582), .B(n4155), .C(n4198), .Y(n4764) );
  INVX1 U1521 ( .A(N3998), .Y(n7582) );
  OAI21X1 U1522 ( .A(n7583), .B(n4155), .C(n4198), .Y(n4763) );
  INVX1 U1523 ( .A(N3995), .Y(n7583) );
  OAI21X1 U1524 ( .A(n7584), .B(n4155), .C(n4198), .Y(n4762) );
  INVX1 U1525 ( .A(N3992), .Y(n7584) );
  OAI21X1 U1526 ( .A(n7585), .B(n4155), .C(n4198), .Y(n4761) );
  NAND2X1 U1527 ( .A(n4168), .B(n4155), .Y(n4198) );
  INVX1 U1528 ( .A(n4199), .Y(n4155) );
  NAND3X1 U1529 ( .A(n3816), .B(n3815), .C(n4170), .Y(n4199) );
  INVX1 U1530 ( .A(n4187), .Y(n4170) );
  INVX1 U1531 ( .A(N3989), .Y(n7585) );
  OAI21X1 U1532 ( .A(n7594), .B(n4156), .C(n4200), .Y(n4760) );
  INVX1 U1533 ( .A(N3986), .Y(n7594) );
  OAI21X1 U1534 ( .A(n7595), .B(n4156), .C(n4200), .Y(n4759) );
  INVX1 U1535 ( .A(N3983), .Y(n7595) );
  OAI21X1 U1536 ( .A(n7596), .B(n4156), .C(n4200), .Y(n4758) );
  INVX1 U1537 ( .A(N3980), .Y(n7596) );
  OAI21X1 U1538 ( .A(n7597), .B(n4156), .C(n4200), .Y(n4757) );
  INVX1 U1539 ( .A(N3977), .Y(n7597) );
  OAI21X1 U1540 ( .A(n7598), .B(n4156), .C(n4200), .Y(n4756) );
  INVX1 U1541 ( .A(N3974), .Y(n7598) );
  OAI21X1 U1542 ( .A(n7599), .B(n4156), .C(n4200), .Y(n4755) );
  INVX1 U1543 ( .A(N3971), .Y(n7599) );
  OAI21X1 U1544 ( .A(n7600), .B(n4156), .C(n4200), .Y(n4754) );
  INVX1 U1545 ( .A(N3968), .Y(n7600) );
  OAI21X1 U1546 ( .A(n7601), .B(n4156), .C(n4200), .Y(n4753) );
  NAND2X1 U1547 ( .A(n4168), .B(n4156), .Y(n4200) );
  NOR2X1 U1548 ( .A(n4187), .B(n3826), .Y(n4156) );
  INVX1 U1549 ( .A(N3965), .Y(n7601) );
  OAI21X1 U1550 ( .A(n7610), .B(n4157), .C(n4201), .Y(n4752) );
  INVX1 U1551 ( .A(N3962), .Y(n7610) );
  OAI21X1 U1552 ( .A(n7611), .B(n4157), .C(n4201), .Y(n4751) );
  INVX1 U1553 ( .A(N3959), .Y(n7611) );
  OAI21X1 U1554 ( .A(n7612), .B(n4157), .C(n4201), .Y(n4750) );
  INVX1 U1555 ( .A(N3956), .Y(n7612) );
  OAI21X1 U1556 ( .A(n7613), .B(n4157), .C(n4201), .Y(n4749) );
  INVX1 U1557 ( .A(N3953), .Y(n7613) );
  OAI21X1 U1558 ( .A(n7614), .B(n4157), .C(n4201), .Y(n4748) );
  INVX1 U1559 ( .A(N3950), .Y(n7614) );
  OAI21X1 U1560 ( .A(n7615), .B(n4157), .C(n4201), .Y(n4747) );
  INVX1 U1561 ( .A(N3947), .Y(n7615) );
  OAI21X1 U1562 ( .A(n7616), .B(n4157), .C(n4201), .Y(n4746) );
  INVX1 U1563 ( .A(N3944), .Y(n7616) );
  OAI21X1 U1564 ( .A(n7617), .B(n4157), .C(n4201), .Y(n4745) );
  NAND2X1 U1565 ( .A(n4168), .B(n4157), .Y(n4201) );
  NOR2X1 U1566 ( .A(n4187), .B(n3840), .Y(n4157) );
  INVX1 U1567 ( .A(N3941), .Y(n7617) );
  OAI21X1 U1568 ( .A(n7626), .B(n4158), .C(n4202), .Y(n4744) );
  INVX1 U1569 ( .A(N3938), .Y(n7626) );
  OAI21X1 U1570 ( .A(n7627), .B(n4158), .C(n4202), .Y(n4743) );
  INVX1 U1571 ( .A(N3935), .Y(n7627) );
  OAI21X1 U1572 ( .A(n7628), .B(n4158), .C(n4202), .Y(n4742) );
  INVX1 U1573 ( .A(N3932), .Y(n7628) );
  OAI21X1 U1574 ( .A(n7629), .B(n4158), .C(n4202), .Y(n4741) );
  INVX1 U1575 ( .A(N3929), .Y(n7629) );
  OAI21X1 U1576 ( .A(n7630), .B(n4158), .C(n4202), .Y(n4740) );
  INVX1 U1577 ( .A(N3926), .Y(n7630) );
  OAI21X1 U1578 ( .A(n7631), .B(n4158), .C(n4202), .Y(n4739) );
  INVX1 U1579 ( .A(N3923), .Y(n7631) );
  OAI21X1 U1580 ( .A(n7632), .B(n4158), .C(n4202), .Y(n4738) );
  INVX1 U1581 ( .A(N3920), .Y(n7632) );
  OAI21X1 U1582 ( .A(n7633), .B(n4158), .C(n4202), .Y(n4737) );
  NAND2X1 U1583 ( .A(n4168), .B(n4158), .Y(n4202) );
  NOR2X1 U1584 ( .A(n4187), .B(n3860), .Y(n4158) );
  INVX1 U1585 ( .A(N3917), .Y(n7633) );
  OAI21X1 U1586 ( .A(n7642), .B(n4159), .C(n4203), .Y(n4736) );
  INVX1 U1587 ( .A(N3914), .Y(n7642) );
  OAI21X1 U1588 ( .A(n7643), .B(n4159), .C(n4203), .Y(n4735) );
  INVX1 U1589 ( .A(N3911), .Y(n7643) );
  OAI21X1 U1590 ( .A(n7644), .B(n4159), .C(n4203), .Y(n4734) );
  INVX1 U1591 ( .A(N3908), .Y(n7644) );
  OAI21X1 U1592 ( .A(n7645), .B(n4159), .C(n4203), .Y(n4733) );
  INVX1 U1593 ( .A(N3905), .Y(n7645) );
  OAI21X1 U1594 ( .A(n7646), .B(n4159), .C(n4203), .Y(n4732) );
  INVX1 U1595 ( .A(N3902), .Y(n7646) );
  OAI21X1 U1596 ( .A(n7647), .B(n4159), .C(n4203), .Y(n4731) );
  INVX1 U1597 ( .A(N3899), .Y(n7647) );
  OAI21X1 U1598 ( .A(n7648), .B(n4159), .C(n4203), .Y(n4730) );
  INVX1 U1599 ( .A(N3896), .Y(n7648) );
  OAI21X1 U1600 ( .A(n7649), .B(n4159), .C(n4203), .Y(n4729) );
  NAND2X1 U1601 ( .A(n4168), .B(n4159), .Y(n4203) );
  NOR2X1 U1602 ( .A(n4187), .B(n4204), .Y(n4159) );
  INVX1 U1603 ( .A(N3893), .Y(n7649) );
  OAI21X1 U1604 ( .A(n7658), .B(n4160), .C(n4205), .Y(n4728) );
  INVX1 U1605 ( .A(N3890), .Y(n7658) );
  OAI21X1 U1606 ( .A(n7659), .B(n4160), .C(n4205), .Y(n4727) );
  INVX1 U1607 ( .A(N3887), .Y(n7659) );
  OAI21X1 U1608 ( .A(n7660), .B(n4160), .C(n4205), .Y(n4726) );
  INVX1 U1609 ( .A(N3884), .Y(n7660) );
  OAI21X1 U1610 ( .A(n7661), .B(n4160), .C(n4205), .Y(n4725) );
  INVX1 U1611 ( .A(N3881), .Y(n7661) );
  OAI21X1 U1612 ( .A(n7662), .B(n4160), .C(n4205), .Y(n4724) );
  INVX1 U1613 ( .A(N3878), .Y(n7662) );
  OAI21X1 U1614 ( .A(n7663), .B(n4160), .C(n4205), .Y(n4723) );
  INVX1 U1615 ( .A(N3875), .Y(n7663) );
  OAI21X1 U1616 ( .A(n7664), .B(n4160), .C(n4205), .Y(n4722) );
  INVX1 U1617 ( .A(N3872), .Y(n7664) );
  OAI21X1 U1618 ( .A(n7665), .B(n4160), .C(n4205), .Y(n4721) );
  NAND2X1 U1619 ( .A(n4168), .B(n4160), .Y(n4205) );
  NOR2X1 U1620 ( .A(n4187), .B(n3890), .Y(n4160) );
  INVX1 U1621 ( .A(N3869), .Y(n7665) );
  OAI21X1 U1622 ( .A(n7674), .B(n4161), .C(n4206), .Y(n4720) );
  INVX1 U1623 ( .A(N3866), .Y(n7674) );
  OAI21X1 U1624 ( .A(n7675), .B(n4161), .C(n4206), .Y(n4719) );
  INVX1 U1625 ( .A(N3863), .Y(n7675) );
  OAI21X1 U1626 ( .A(n7676), .B(n4161), .C(n4206), .Y(n4718) );
  INVX1 U1627 ( .A(N3860), .Y(n7676) );
  OAI21X1 U1628 ( .A(n7677), .B(n4161), .C(n4206), .Y(n4717) );
  INVX1 U1629 ( .A(N3857), .Y(n7677) );
  OAI21X1 U1630 ( .A(n7678), .B(n4161), .C(n4206), .Y(n4716) );
  INVX1 U1631 ( .A(N3854), .Y(n7678) );
  OAI21X1 U1632 ( .A(n7679), .B(n4161), .C(n4206), .Y(n4715) );
  INVX1 U1633 ( .A(N3851), .Y(n7679) );
  OAI21X1 U1634 ( .A(n7680), .B(n4161), .C(n4206), .Y(n4714) );
  INVX1 U1635 ( .A(N3848), .Y(n7680) );
  OAI21X1 U1636 ( .A(n7681), .B(n4161), .C(n4206), .Y(n4713) );
  NAND2X1 U1637 ( .A(n4168), .B(n4161), .Y(n4206) );
  NOR2X1 U1638 ( .A(n4187), .B(n3902), .Y(n4161) );
  INVX1 U1639 ( .A(N3845), .Y(n7681) );
  OAI21X1 U1640 ( .A(n7322), .B(n4162), .C(n4207), .Y(n4712) );
  INVX1 U1641 ( .A(N3842), .Y(n7322) );
  OAI21X1 U1642 ( .A(n7323), .B(n4162), .C(n4207), .Y(n4711) );
  INVX1 U1643 ( .A(N3839), .Y(n7323) );
  OAI21X1 U1644 ( .A(n7324), .B(n4162), .C(n4207), .Y(n4710) );
  INVX1 U1645 ( .A(N3836), .Y(n7324) );
  OAI21X1 U1646 ( .A(n7325), .B(n4162), .C(n4207), .Y(n4709) );
  INVX1 U1647 ( .A(N3833), .Y(n7325) );
  OAI21X1 U1648 ( .A(n7326), .B(n4162), .C(n4207), .Y(n4708) );
  INVX1 U1649 ( .A(N3830), .Y(n7326) );
  OAI21X1 U1650 ( .A(n7327), .B(n4162), .C(n4207), .Y(n4707) );
  INVX1 U1651 ( .A(N3827), .Y(n7327) );
  OAI21X1 U1652 ( .A(n7328), .B(n4162), .C(n4207), .Y(n4706) );
  INVX1 U1653 ( .A(N3824), .Y(n7328) );
  OAI21X1 U1654 ( .A(n7329), .B(n4162), .C(n4207), .Y(n4705) );
  NAND2X1 U1655 ( .A(n4168), .B(n4162), .Y(n4207) );
  NOR2X1 U1656 ( .A(n4187), .B(n3912), .Y(n4162) );
  INVX1 U1657 ( .A(N3821), .Y(n7329) );
  OAI21X1 U1658 ( .A(n7306), .B(n4163), .C(n4208), .Y(n4704) );
  INVX1 U1659 ( .A(N3818), .Y(n7306) );
  OAI21X1 U1660 ( .A(n7307), .B(n4163), .C(n4208), .Y(n4703) );
  INVX1 U1661 ( .A(N3815), .Y(n7307) );
  OAI21X1 U1662 ( .A(n7308), .B(n4163), .C(n4208), .Y(n4702) );
  INVX1 U1663 ( .A(N3812), .Y(n7308) );
  OAI21X1 U1664 ( .A(n7309), .B(n4163), .C(n4208), .Y(n4701) );
  INVX1 U1665 ( .A(N3809), .Y(n7309) );
  OAI21X1 U1666 ( .A(n7310), .B(n4163), .C(n4208), .Y(n4700) );
  INVX1 U1667 ( .A(N3806), .Y(n7310) );
  OAI21X1 U1668 ( .A(n7311), .B(n4163), .C(n4208), .Y(n4699) );
  INVX1 U1669 ( .A(N3803), .Y(n7311) );
  OAI21X1 U1670 ( .A(n7312), .B(n4163), .C(n4208), .Y(n4698) );
  INVX1 U1671 ( .A(N3800), .Y(n7312) );
  OAI21X1 U1672 ( .A(n7313), .B(n4163), .C(n4208), .Y(n4697) );
  NAND2X1 U1673 ( .A(n4168), .B(n4163), .Y(n4208) );
  NOR2X1 U1674 ( .A(n4187), .B(n3925), .Y(n4163) );
  INVX1 U1675 ( .A(N3797), .Y(n7313) );
  OAI21X1 U1676 ( .A(n7690), .B(n4164), .C(n4209), .Y(n4696) );
  INVX1 U1677 ( .A(N3794), .Y(n7690) );
  OAI21X1 U1678 ( .A(n7691), .B(n4164), .C(n4209), .Y(n4695) );
  INVX1 U1679 ( .A(N3791), .Y(n7691) );
  OAI21X1 U1680 ( .A(n7692), .B(n4164), .C(n4209), .Y(n4694) );
  INVX1 U1681 ( .A(N3788), .Y(n7692) );
  OAI21X1 U1682 ( .A(n7693), .B(n4164), .C(n4209), .Y(n4693) );
  INVX1 U1683 ( .A(N3785), .Y(n7693) );
  OAI21X1 U1684 ( .A(n7694), .B(n4164), .C(n4209), .Y(n4692) );
  INVX1 U1685 ( .A(N3782), .Y(n7694) );
  OAI21X1 U1686 ( .A(n7695), .B(n4164), .C(n4209), .Y(n4691) );
  INVX1 U1687 ( .A(N3779), .Y(n7695) );
  OAI21X1 U1688 ( .A(n7696), .B(n4164), .C(n4209), .Y(n4690) );
  INVX1 U1689 ( .A(N3776), .Y(n7696) );
  OAI21X1 U1690 ( .A(n7697), .B(n4164), .C(n4209), .Y(n4689) );
  NAND2X1 U1691 ( .A(n4168), .B(n4164), .Y(n4209) );
  NOR2X1 U1692 ( .A(n4187), .B(n3941), .Y(n4164) );
  OAI21X1 U1693 ( .A(n4168), .B(n4210), .C(rst_b), .Y(n4187) );
  NOR2X1 U1694 ( .A(n4166), .B(n4211), .Y(n4210) );
  NAND2X1 U1695 ( .A(n3490), .B(n3853), .Y(n4211) );
  NAND2X1 U1696 ( .A(dWriteReg[1]), .B(n3945), .Y(n4166) );
  INVX1 U1697 ( .A(n4212), .Y(n4168) );
  NAND3X1 U1698 ( .A(n3490), .B(n3853), .C(n4213), .Y(n4212) );
  AOI21X1 U1699 ( .A(n4214), .B(n3944), .C(n3945), .Y(n4213) );
  NOR3X1 U1700 ( .A(dWriteReg[2]), .B(dWriteReg[3]), .C(dWriteReg[0]), .Y(
        n3945) );
  INVX1 U1701 ( .A(N3773), .Y(n7697) );
  OAI21X1 U1702 ( .A(n7281), .B(n3558), .C(n3559), .Y(n4681) );
  NAND3X1 U1703 ( .A(n3558), .B(n4215), .C(n4216), .Y(n3559) );
  NOR2X1 U1704 ( .A(n4217), .B(n4218), .Y(n4216) );
  NAND2X1 U1705 ( .A(n4219), .B(n4220), .Y(n4218) );
  INVX1 U1706 ( .A(N4496), .Y(n7281) );
  OR2X1 U1707 ( .A(n4221), .B(n4222), .Y(n4680) );
  OAI22X1 U1708 ( .A(n7280), .B(n3558), .C(n4215), .D(n4223), .Y(n4222) );
  INVX1 U1709 ( .A(N4495), .Y(n7280) );
  OAI21X1 U1710 ( .A(n4224), .B(n4225), .C(n4226), .Y(n4221) );
  OAI21X1 U1711 ( .A(n3558), .B(n4227), .C(n4226), .Y(n4679) );
  INVX1 U1712 ( .A(dy[1]), .Y(n4227) );
  OR2X1 U1713 ( .A(n4228), .B(n4229), .Y(n4678) );
  OAI22X1 U1714 ( .A(n7279), .B(n3558), .C(n4224), .D(n4223), .Y(n4229) );
  INVX1 U1715 ( .A(n4217), .Y(n4224) );
  NOR2X1 U1716 ( .A(n4230), .B(n4231), .Y(n4217) );
  NAND3X1 U1717 ( .A(n4232), .B(\regY[6][1] ), .C(\regY[6][4] ), .Y(n4231) );
  NAND3X1 U1718 ( .A(\regY[6][6] ), .B(n4233), .C(\regY[6][3] ), .Y(n4230) );
  INVX1 U1719 ( .A(N4501), .Y(n7279) );
  OAI21X1 U1720 ( .A(n4225), .B(n4215), .C(n4226), .Y(n4228) );
  OAI21X1 U1721 ( .A(n4234), .B(n4235), .C(n3558), .Y(n4226) );
  INVX1 U1722 ( .A(n4219), .Y(n4235) );
  NAND3X1 U1723 ( .A(n4236), .B(n4237), .C(n4232), .Y(n4215) );
  INVX1 U1724 ( .A(n4238), .Y(n4232) );
  NAND3X1 U1725 ( .A(n4239), .B(n4240), .C(n4241), .Y(n4238) );
  OAI21X1 U1726 ( .A(n3558), .B(n4242), .C(n4243), .Y(n4677) );
  INVX1 U1727 ( .A(n4244), .Y(n4243) );
  OAI22X1 U1728 ( .A(n4219), .B(n4225), .C(n4220), .D(n4223), .Y(n4244) );
  NAND2X1 U1729 ( .A(n3558), .B(OPMode[0]), .Y(n4223) );
  INVX1 U1730 ( .A(n4234), .Y(n4220) );
  NOR2X1 U1731 ( .A(n4245), .B(n4246), .Y(n4234) );
  NAND3X1 U1732 ( .A(\regY[6][5] ), .B(\regY[6][3] ), .C(n4247), .Y(n4246) );
  NAND3X1 U1733 ( .A(n4237), .B(n4248), .C(n4249), .Y(n4245) );
  NOR2X1 U1734 ( .A(\regY[6][7] ), .B(\regY[6][6] ), .Y(n4249) );
  NAND2X1 U1735 ( .A(n3558), .B(n4250), .Y(n4225) );
  NAND3X1 U1736 ( .A(n4247), .B(n4236), .C(n4251), .Y(n4219) );
  NOR2X1 U1737 ( .A(n4237), .B(n4240), .Y(n4251) );
  INVX1 U1738 ( .A(n4252), .Y(n4236) );
  NAND3X1 U1739 ( .A(n4253), .B(n4248), .C(n4254), .Y(n4252) );
  NOR2X1 U1740 ( .A(\regY[6][6] ), .B(\regY[6][5] ), .Y(n4254) );
  NOR2X1 U1741 ( .A(n4241), .B(n4239), .Y(n4247) );
  INVX1 U1742 ( .A(n4255), .Y(n3558) );
  NAND3X1 U1743 ( .A(n4256), .B(n4257), .C(n3936), .Y(n4255) );
  OAI21X1 U1744 ( .A(n7713), .B(n4258), .C(n4259), .Y(n4676) );
  INVX1 U1745 ( .A(N4418), .Y(n7713) );
  OAI21X1 U1746 ( .A(n7712), .B(n4258), .C(n4259), .Y(n4675) );
  INVX1 U1747 ( .A(N4415), .Y(n7712) );
  OAI21X1 U1748 ( .A(n7711), .B(n4258), .C(n4259), .Y(n4674) );
  INVX1 U1749 ( .A(N4412), .Y(n7711) );
  OAI21X1 U1750 ( .A(n7710), .B(n4258), .C(n4259), .Y(n4673) );
  INVX1 U1751 ( .A(N4409), .Y(n7710) );
  OAI21X1 U1752 ( .A(n7709), .B(n4258), .C(n4259), .Y(n4672) );
  INVX1 U1753 ( .A(N4406), .Y(n7709) );
  OAI21X1 U1754 ( .A(n7708), .B(n4258), .C(n4259), .Y(n4671) );
  INVX1 U1755 ( .A(N4403), .Y(n7708) );
  OAI21X1 U1756 ( .A(n7707), .B(n4258), .C(n4259), .Y(n4670) );
  INVX1 U1757 ( .A(N4400), .Y(n7707) );
  OAI21X1 U1758 ( .A(n7706), .B(n4258), .C(n4259), .Y(n4669) );
  NAND2X1 U1759 ( .A(n4258), .B(n3484), .Y(n4259) );
  INVX1 U1760 ( .A(N4397), .Y(n7706) );
  OAI21X1 U1761 ( .A(n7705), .B(n4258), .C(n4260), .Y(n4668) );
  AOI22X1 U1762 ( .A(N2569), .B(n4261), .C(N2561), .D(n4262), .Y(n4260) );
  INVX1 U1763 ( .A(N4417), .Y(n7705) );
  OAI21X1 U1764 ( .A(n7704), .B(n4258), .C(n4263), .Y(n4667) );
  AOI22X1 U1765 ( .A(N2570), .B(n4261), .C(N2562), .D(n4262), .Y(n4263) );
  INVX1 U1766 ( .A(N4414), .Y(n7704) );
  OAI21X1 U1767 ( .A(n7703), .B(n4258), .C(n4264), .Y(n4666) );
  AOI22X1 U1768 ( .A(N2571), .B(n4261), .C(N2563), .D(n4262), .Y(n4264) );
  INVX1 U1769 ( .A(N4411), .Y(n7703) );
  OAI21X1 U1770 ( .A(n7702), .B(n4258), .C(n4265), .Y(n4665) );
  AOI22X1 U1771 ( .A(N2572), .B(n4261), .C(N2564), .D(n4262), .Y(n4265) );
  INVX1 U1772 ( .A(N4408), .Y(n7702) );
  OAI21X1 U1773 ( .A(n7701), .B(n4258), .C(n4266), .Y(n4664) );
  AOI22X1 U1774 ( .A(N2573), .B(n4261), .C(N2565), .D(n4262), .Y(n4266) );
  INVX1 U1775 ( .A(N4405), .Y(n7701) );
  OAI21X1 U1776 ( .A(n7700), .B(n4258), .C(n4267), .Y(n4663) );
  AOI22X1 U1777 ( .A(N2574), .B(n4261), .C(N2566), .D(n4262), .Y(n4267) );
  INVX1 U1778 ( .A(N4402), .Y(n7700) );
  OAI21X1 U1779 ( .A(n7699), .B(n4258), .C(n4268), .Y(n4662) );
  AOI22X1 U1780 ( .A(N2575), .B(n4261), .C(N2567), .D(n4262), .Y(n4268) );
  INVX1 U1781 ( .A(N4399), .Y(n7699) );
  OAI21X1 U1782 ( .A(n7698), .B(n4258), .C(n4269), .Y(n4661) );
  AOI22X1 U1783 ( .A(N2576), .B(n4261), .C(N2568), .D(n4262), .Y(n4269) );
  INVX1 U1784 ( .A(n4270), .Y(n4262) );
  NAND3X1 U1785 ( .A(n3707), .B(n4128), .C(n4258), .Y(n4270) );
  INVX1 U1786 ( .A(n4271), .Y(n4261) );
  OAI21X1 U1787 ( .A(n4080), .B(n4272), .C(n4258), .Y(n4271) );
  AND2X1 U1788 ( .A(n3936), .B(n4273), .Y(n4258) );
  INVX1 U1789 ( .A(N4396), .Y(n7698) );
  OAI21X1 U1790 ( .A(n4274), .B(n4275), .C(n4276), .Y(n4660) );
  NAND2X1 U1791 ( .A(N2048), .B(n4277), .Y(n4276) );
  OAI21X1 U1792 ( .A(n4274), .B(n4278), .C(n4279), .Y(n4659) );
  NAND2X1 U1793 ( .A(N2049), .B(n4277), .Y(n4279) );
  OAI21X1 U1794 ( .A(n4274), .B(n4280), .C(n4281), .Y(n4658) );
  NAND2X1 U1795 ( .A(N2050), .B(n4277), .Y(n4281) );
  OAI21X1 U1796 ( .A(n4274), .B(n4282), .C(n4283), .Y(n4657) );
  NAND2X1 U1797 ( .A(N2051), .B(n4277), .Y(n4283) );
  OAI21X1 U1798 ( .A(n4274), .B(n4284), .C(n4285), .Y(n4656) );
  NAND2X1 U1799 ( .A(N2052), .B(n4277), .Y(n4285) );
  OAI21X1 U1800 ( .A(n4274), .B(n4286), .C(n4287), .Y(n4655) );
  NAND2X1 U1801 ( .A(N2053), .B(n4277), .Y(n4287) );
  OAI21X1 U1802 ( .A(n4274), .B(n4288), .C(n4289), .Y(n4654) );
  NAND2X1 U1803 ( .A(N2054), .B(n4277), .Y(n4289) );
  OAI21X1 U1804 ( .A(n4274), .B(n4290), .C(n4291), .Y(n4653) );
  NAND2X1 U1805 ( .A(N2055), .B(n4277), .Y(n4291) );
  NOR2X1 U1806 ( .A(n4292), .B(n3548), .Y(n4277) );
  NOR2X1 U1807 ( .A(n4292), .B(n4293), .Y(n4274) );
  MUX2X1 U1808 ( .B(n4294), .A(n4295), .S(n4296), .Y(n4652) );
  NOR2X1 U1809 ( .A(n4297), .B(n3850), .Y(n4296) );
  OAI22X1 U1810 ( .A(n4080), .B(n4298), .C(n4299), .D(n4300), .Y(n4295) );
  NAND2X1 U1811 ( .A(n4301), .B(N2880), .Y(n4300) );
  OAI22X1 U1812 ( .A(n4302), .B(n4303), .C(n4304), .D(n4305), .Y(n4299) );
  NAND2X1 U1813 ( .A(n4306), .B(n4307), .Y(n4305) );
  OAI21X1 U1814 ( .A(n4308), .B(n4309), .C(n4310), .Y(n4307) );
  OAI21X1 U1815 ( .A(n4311), .B(n4312), .C(n4313), .Y(n4309) );
  NAND3X1 U1816 ( .A(n4314), .B(n4315), .C(n4316), .Y(n4313) );
  INVX1 U1817 ( .A(n4317), .Y(n4311) );
  MUX2X1 U1818 ( .B(n4318), .A(n4319), .S(n4320), .Y(n4308) );
  AND2X1 U1819 ( .A(n4321), .B(n4322), .Y(n4319) );
  AOI22X1 U1820 ( .A(n4323), .B(n4324), .C(n4325), .D(n4326), .Y(n4322) );
  AOI22X1 U1821 ( .A(n4327), .B(n4328), .C(n4329), .D(n4316), .Y(n4321) );
  AOI21X1 U1822 ( .A(n4324), .B(n4330), .C(n4331), .Y(n4318) );
  OAI21X1 U1823 ( .A(n4332), .B(n4333), .C(n4334), .Y(n4331) );
  NAND3X1 U1824 ( .A(n4312), .B(n4335), .C(n4326), .Y(n4334) );
  INVX1 U1825 ( .A(n4336), .Y(n4332) );
  MUX2X1 U1826 ( .B(n4337), .A(n4338), .S(n4339), .Y(n4306) );
  MUX2X1 U1827 ( .B(n4340), .A(n4341), .S(n4320), .Y(n4338) );
  AND2X1 U1828 ( .A(n4342), .B(n4343), .Y(n4341) );
  AOI22X1 U1829 ( .A(n4344), .B(n4316), .C(n4345), .D(n4326), .Y(n4343) );
  AOI22X1 U1830 ( .A(n4346), .B(n4324), .C(n4347), .D(n4328), .Y(n4342) );
  NOR2X1 U1831 ( .A(n4348), .B(n4349), .Y(n4340) );
  OAI22X1 U1832 ( .A(n4350), .B(n4351), .C(n4352), .D(n4333), .Y(n4349) );
  INVX1 U1833 ( .A(n4353), .Y(n4352) );
  OAI21X1 U1834 ( .A(n4354), .B(n4355), .C(n4356), .Y(n4348) );
  NAND3X1 U1835 ( .A(n4357), .B(n4358), .C(n4326), .Y(n4356) );
  INVX1 U1836 ( .A(n4359), .Y(n4354) );
  NOR2X1 U1837 ( .A(n4310), .B(n4360), .Y(n4337) );
  OAI21X1 U1838 ( .A(n4361), .B(n4362), .C(n4315), .Y(n4360) );
  OAI22X1 U1839 ( .A(n4363), .B(n4333), .C(n4364), .D(n4351), .Y(n4362) );
  AND2X1 U1840 ( .A(n4365), .B(n4326), .Y(n4361) );
  OAI21X1 U1841 ( .A(n4366), .B(n4367), .C(n4368), .Y(n4304) );
  OAI21X1 U1842 ( .A(n4369), .B(n4370), .C(n4371), .Y(n4368) );
  INVX1 U1843 ( .A(n4372), .Y(n4371) );
  OAI22X1 U1844 ( .A(n4373), .B(n4333), .C(n4374), .D(n4351), .Y(n4370) );
  INVX1 U1845 ( .A(n4375), .Y(n4369) );
  AOI22X1 U1846 ( .A(n4376), .B(n4326), .C(n4377), .D(n4316), .Y(n4375) );
  OAI21X1 U1847 ( .A(n4378), .B(n4379), .C(n4380), .Y(n4367) );
  OAI21X1 U1848 ( .A(n4381), .B(n4382), .C(n4383), .Y(n4380) );
  OAI21X1 U1849 ( .A(n4312), .B(n4384), .C(n4357), .Y(n4383) );
  OAI21X1 U1850 ( .A(n4355), .B(n4385), .C(n4386), .Y(n4382) );
  OAI21X1 U1851 ( .A(\regZ[24][0] ), .B(n4387), .C(n4339), .Y(n4386) );
  INVX1 U1852 ( .A(n4312), .Y(n4339) );
  INVX1 U1853 ( .A(n4384), .Y(n4387) );
  MUX2X1 U1854 ( .B(n4388), .A(n4389), .S(n4320), .Y(n4384) );
  NAND2X1 U1855 ( .A(n4390), .B(n4391), .Y(n4389) );
  AOI22X1 U1856 ( .A(\regZ[17][0] ), .B(n4326), .C(\regZ[23][0] ), .D(n4316), 
        .Y(n4391) );
  AOI22X1 U1857 ( .A(\regZ[19][0] ), .B(n4324), .C(\regZ[21][0] ), .D(n4328), 
        .Y(n4390) );
  NAND2X1 U1858 ( .A(n4392), .B(n4393), .Y(n4388) );
  AOI22X1 U1859 ( .A(n4394), .B(\regZ[16][0] ), .C(\regZ[22][0] ), .D(n4316), 
        .Y(n4393) );
  NOR2X1 U1860 ( .A(n4395), .B(n4310), .Y(n4394) );
  AOI22X1 U1861 ( .A(\regZ[18][0] ), .B(n4324), .C(\regZ[20][0] ), .D(n4328), 
        .Y(n4392) );
  MUX2X1 U1862 ( .B(\regZ[14][0] ), .A(\regZ[15][0] ), .S(n4320), .Y(n4385) );
  MUX2X1 U1863 ( .B(n4396), .A(n4397), .S(n4320), .Y(n4381) );
  AOI21X1 U1864 ( .A(\regZ[13][0] ), .B(n4328), .C(n4398), .Y(n4397) );
  OAI22X1 U1865 ( .A(n4351), .B(n4399), .C(n4395), .D(n4400), .Y(n4398) );
  AOI22X1 U1866 ( .A(\regZ[10][0] ), .B(n4324), .C(\regZ[12][0] ), .D(n4328), 
        .Y(n4396) );
  NAND2X1 U1867 ( .A(n4312), .B(n4315), .Y(n4379) );
  MUX2X1 U1868 ( .B(n4401), .A(n4402), .S(n4310), .Y(n4378) );
  INVX1 U1869 ( .A(n4357), .Y(n4310) );
  NOR2X1 U1870 ( .A(n4395), .B(n4403), .Y(n4402) );
  OAI21X1 U1871 ( .A(n4333), .B(n4404), .C(n4405), .Y(n4401) );
  AOI22X1 U1872 ( .A(\regZ[0][0] ), .B(n4326), .C(\regZ[2][0] ), .D(n4324), 
        .Y(n4405) );
  INVX1 U1873 ( .A(\regZ[4][0] ), .Y(n4404) );
  AOI21X1 U1874 ( .A(n4406), .B(n4407), .C(n4372), .Y(n4366) );
  NAND3X1 U1875 ( .A(n4357), .B(n4312), .C(n4320), .Y(n4372) );
  INVX1 U1876 ( .A(n4315), .Y(n4320) );
  OAI21X1 U1877 ( .A(n4408), .B(dx[0]), .C(n4409), .Y(n4315) );
  XOR2X1 U1878 ( .A(n4410), .B(n4411), .Y(n4312) );
  XOR2X1 U1879 ( .A(n4242), .B(n4412), .Y(n4411) );
  XOR2X1 U1880 ( .A(n4413), .B(n4414), .Y(n4410) );
  NOR2X1 U1881 ( .A(n4415), .B(n4416), .Y(n4414) );
  OAI21X1 U1882 ( .A(n4417), .B(n4418), .C(n4419), .Y(n4413) );
  OAI21X1 U1883 ( .A(n4420), .B(n4421), .C(dx[1]), .Y(n4419) );
  XOR2X1 U1884 ( .A(n4422), .B(n4421), .Y(n4357) );
  XOR2X1 U1885 ( .A(n4242), .B(n4420), .Y(n4422) );
  INVX1 U1886 ( .A(n4418), .Y(n4420) );
  OAI21X1 U1887 ( .A(n4423), .B(n4424), .C(n4425), .Y(n4418) );
  OAI21X1 U1888 ( .A(n4426), .B(n4427), .C(n4242), .Y(n4425) );
  INVX1 U1889 ( .A(n4424), .Y(n4427) );
  AOI22X1 U1890 ( .A(\regZ[1][0] ), .B(n4326), .C(\regZ[7][0] ), .D(n4316), 
        .Y(n4407) );
  INVX1 U1891 ( .A(n4355), .Y(n4316) );
  NAND2X1 U1892 ( .A(n4428), .B(n4429), .Y(n4355) );
  INVX1 U1893 ( .A(n4395), .Y(n4326) );
  NAND2X1 U1894 ( .A(n4430), .B(n4431), .Y(n4395) );
  AOI22X1 U1895 ( .A(\regZ[3][0] ), .B(n4324), .C(\regZ[5][0] ), .D(n4328), 
        .Y(n4406) );
  INVX1 U1896 ( .A(n4333), .Y(n4328) );
  NAND2X1 U1897 ( .A(n4429), .B(n4431), .Y(n4333) );
  INVX1 U1898 ( .A(n4430), .Y(n4429) );
  INVX1 U1899 ( .A(n4351), .Y(n4324) );
  NAND2X1 U1900 ( .A(n4430), .B(n4428), .Y(n4351) );
  INVX1 U1901 ( .A(n4431), .Y(n4428) );
  XOR2X1 U1902 ( .A(n4432), .B(n4433), .Y(n4431) );
  XOR2X1 U1903 ( .A(n4242), .B(n4434), .Y(n4432) );
  XOR2X1 U1904 ( .A(n4435), .B(n4426), .Y(n4430) );
  INVX1 U1905 ( .A(n4423), .Y(n4426) );
  OAI21X1 U1906 ( .A(n4436), .B(n4409), .C(n4437), .Y(n4423) );
  OAI21X1 U1907 ( .A(n4434), .B(n4433), .C(dx[1]), .Y(n4437) );
  INVX1 U1908 ( .A(n4409), .Y(n4434) );
  NAND2X1 U1909 ( .A(n4408), .B(dx[0]), .Y(n4409) );
  XOR2X1 U1910 ( .A(n4424), .B(dx[1]), .Y(n4435) );
  OAI21X1 U1911 ( .A(n4373), .B(n4438), .C(n4439), .Y(n4303) );
  AOI22X1 U1912 ( .A(n4440), .B(n4441), .C(n3586), .D(n4442), .Y(n4439) );
  NAND3X1 U1913 ( .A(n4443), .B(n4444), .C(n4445), .Y(n4442) );
  NOR2X1 U1914 ( .A(n4446), .B(n4447), .Y(n4445) );
  OAI21X1 U1915 ( .A(n4350), .B(n3652), .C(n4448), .Y(n4447) );
  MUX2X1 U1916 ( .B(n4449), .A(n4317), .S(n3585), .Y(n4448) );
  NAND3X1 U1917 ( .A(n4450), .B(n4451), .C(n4452), .Y(n4317) );
  NOR2X1 U1918 ( .A(\regZ[24][1] ), .B(n4453), .Y(n4452) );
  OR2X1 U1919 ( .A(\regZ[24][3] ), .B(\regZ[24][2] ), .Y(n4453) );
  NOR2X1 U1920 ( .A(\regZ[24][7] ), .B(\regZ[24][6] ), .Y(n4451) );
  NOR2X1 U1921 ( .A(\regZ[24][5] ), .B(\regZ[24][4] ), .Y(n4450) );
  AND2X1 U1922 ( .A(n4358), .B(n3583), .Y(n4449) );
  NAND3X1 U1923 ( .A(n4454), .B(n4455), .C(n4456), .Y(n4358) );
  NOR2X1 U1924 ( .A(\regZ[16][1] ), .B(n4457), .Y(n4456) );
  OR2X1 U1925 ( .A(\regZ[16][3] ), .B(\regZ[16][2] ), .Y(n4457) );
  NOR2X1 U1926 ( .A(\regZ[16][7] ), .B(\regZ[16][6] ), .Y(n4455) );
  NOR2X1 U1927 ( .A(\regZ[16][5] ), .B(\regZ[16][4] ), .Y(n4454) );
  INVX1 U1928 ( .A(n4458), .Y(n4350) );
  NAND3X1 U1929 ( .A(n4459), .B(n4460), .C(n4461), .Y(n4458) );
  NOR2X1 U1930 ( .A(\regZ[18][1] ), .B(n4462), .Y(n4461) );
  OR2X1 U1931 ( .A(\regZ[18][3] ), .B(\regZ[18][2] ), .Y(n4462) );
  NOR2X1 U1932 ( .A(\regZ[18][7] ), .B(\regZ[18][6] ), .Y(n4460) );
  NOR2X1 U1933 ( .A(\regZ[18][5] ), .B(\regZ[18][4] ), .Y(n4459) );
  INVX1 U1934 ( .A(n4463), .Y(n4446) );
  AOI22X1 U1935 ( .A(n4345), .B(n3924), .C(n4346), .D(n3901), .Y(n4463) );
  NAND3X1 U1936 ( .A(n4464), .B(n4465), .C(n4466), .Y(n4346) );
  NOR2X1 U1937 ( .A(\regZ[19][1] ), .B(n4467), .Y(n4466) );
  OR2X1 U1938 ( .A(\regZ[19][3] ), .B(\regZ[19][2] ), .Y(n4467) );
  NOR2X1 U1939 ( .A(\regZ[19][7] ), .B(\regZ[19][6] ), .Y(n4465) );
  NOR2X1 U1940 ( .A(\regZ[19][5] ), .B(\regZ[19][4] ), .Y(n4464) );
  NAND3X1 U1941 ( .A(n4468), .B(n4469), .C(n4470), .Y(n4345) );
  NOR2X1 U1942 ( .A(\regZ[17][1] ), .B(n4471), .Y(n4470) );
  OR2X1 U1943 ( .A(\regZ[17][3] ), .B(\regZ[17][2] ), .Y(n4471) );
  NOR2X1 U1944 ( .A(\regZ[17][7] ), .B(\regZ[17][6] ), .Y(n4469) );
  NOR2X1 U1945 ( .A(\regZ[17][5] ), .B(\regZ[17][4] ), .Y(n4468) );
  AOI22X1 U1946 ( .A(n3838), .B(n4344), .C(n3865), .D(n4359), .Y(n4444) );
  NAND3X1 U1947 ( .A(n4472), .B(n4473), .C(n4474), .Y(n4359) );
  NOR2X1 U1948 ( .A(\regZ[22][1] ), .B(n4475), .Y(n4474) );
  OR2X1 U1949 ( .A(\regZ[22][3] ), .B(\regZ[22][2] ), .Y(n4475) );
  NOR2X1 U1950 ( .A(\regZ[22][7] ), .B(\regZ[22][6] ), .Y(n4473) );
  NOR2X1 U1951 ( .A(\regZ[22][5] ), .B(\regZ[22][4] ), .Y(n4472) );
  NAND3X1 U1952 ( .A(n4476), .B(n4477), .C(n4478), .Y(n4344) );
  NOR2X1 U1953 ( .A(\regZ[23][1] ), .B(n4479), .Y(n4478) );
  OR2X1 U1954 ( .A(\regZ[23][3] ), .B(\regZ[23][2] ), .Y(n4479) );
  NOR2X1 U1955 ( .A(\regZ[23][7] ), .B(\regZ[23][6] ), .Y(n4477) );
  NOR2X1 U1956 ( .A(\regZ[23][5] ), .B(\regZ[23][4] ), .Y(n4476) );
  AOI22X1 U1957 ( .A(n4480), .B(n4347), .C(n3889), .D(n4353), .Y(n4443) );
  NAND3X1 U1958 ( .A(n4481), .B(n4482), .C(n4483), .Y(n4353) );
  NOR2X1 U1959 ( .A(\regZ[20][1] ), .B(n4484), .Y(n4483) );
  OR2X1 U1960 ( .A(\regZ[20][3] ), .B(\regZ[20][2] ), .Y(n4484) );
  NOR2X1 U1961 ( .A(\regZ[20][7] ), .B(\regZ[20][6] ), .Y(n4482) );
  NOR2X1 U1962 ( .A(\regZ[20][5] ), .B(\regZ[20][4] ), .Y(n4481) );
  NAND3X1 U1963 ( .A(n4485), .B(n4486), .C(n4487), .Y(n4347) );
  NOR2X1 U1964 ( .A(\regZ[21][1] ), .B(n4488), .Y(n4487) );
  OR2X1 U1965 ( .A(\regZ[21][3] ), .B(\regZ[21][2] ), .Y(n4488) );
  NOR2X1 U1966 ( .A(\regZ[21][7] ), .B(\regZ[21][6] ), .Y(n4486) );
  NOR2X1 U1967 ( .A(\regZ[21][5] ), .B(\regZ[21][4] ), .Y(n4485) );
  NOR2X1 U1968 ( .A(n4363), .B(n3631), .Y(n4440) );
  INVX1 U1969 ( .A(n4489), .Y(n4363) );
  NAND3X1 U1970 ( .A(n4490), .B(n4491), .C(n4492), .Y(n4489) );
  NOR2X1 U1971 ( .A(\regZ[4][1] ), .B(n4493), .Y(n4492) );
  OR2X1 U1972 ( .A(\regZ[4][3] ), .B(\regZ[4][2] ), .Y(n4493) );
  NOR2X1 U1973 ( .A(\regZ[4][7] ), .B(\regZ[4][6] ), .Y(n4491) );
  NOR2X1 U1974 ( .A(\regZ[4][5] ), .B(\regZ[4][4] ), .Y(n4490) );
  INVX1 U1975 ( .A(n4494), .Y(n4373) );
  NAND3X1 U1976 ( .A(n4495), .B(n4496), .C(n4497), .Y(n4494) );
  NOR2X1 U1977 ( .A(\regZ[5][1] ), .B(n4498), .Y(n4497) );
  OR2X1 U1978 ( .A(\regZ[5][3] ), .B(\regZ[5][2] ), .Y(n4498) );
  NOR2X1 U1979 ( .A(\regZ[5][7] ), .B(\regZ[5][6] ), .Y(n4496) );
  NOR2X1 U1980 ( .A(\regZ[5][5] ), .B(\regZ[5][4] ), .Y(n4495) );
  OR2X1 U1981 ( .A(n4499), .B(n4500), .Y(n4302) );
  OAI21X1 U1982 ( .A(n4364), .B(n3913), .C(n4501), .Y(n4500) );
  OAI21X1 U1983 ( .A(n4502), .B(n4503), .C(n3585), .Y(n4501) );
  NAND2X1 U1984 ( .A(n4504), .B(n4505), .Y(n4503) );
  AOI22X1 U1985 ( .A(n3889), .B(n4336), .C(n3901), .D(n4323), .Y(n4505) );
  NAND3X1 U1986 ( .A(n4506), .B(n4507), .C(n4508), .Y(n4323) );
  NOR2X1 U1987 ( .A(\regZ[11][1] ), .B(n4509), .Y(n4508) );
  OR2X1 U1988 ( .A(\regZ[11][3] ), .B(\regZ[11][2] ), .Y(n4509) );
  NOR2X1 U1989 ( .A(\regZ[11][7] ), .B(\regZ[11][6] ), .Y(n4507) );
  NOR2X1 U1990 ( .A(\regZ[11][5] ), .B(\regZ[11][4] ), .Y(n4506) );
  NAND3X1 U1991 ( .A(n4510), .B(n4511), .C(n4512), .Y(n4336) );
  NOR2X1 U1992 ( .A(\regZ[12][1] ), .B(n4513), .Y(n4512) );
  OR2X1 U1993 ( .A(\regZ[12][3] ), .B(\regZ[12][2] ), .Y(n4513) );
  NOR2X1 U1994 ( .A(\regZ[12][7] ), .B(\regZ[12][6] ), .Y(n4511) );
  NOR2X1 U1995 ( .A(\regZ[12][5] ), .B(\regZ[12][4] ), .Y(n4510) );
  AOI22X1 U1996 ( .A(n3924), .B(n4325), .C(n4514), .D(n4330), .Y(n4504) );
  NAND3X1 U1997 ( .A(n4515), .B(n4516), .C(n4517), .Y(n4330) );
  NOR2X1 U1998 ( .A(\regZ[10][1] ), .B(n4518), .Y(n4517) );
  OR2X1 U1999 ( .A(\regZ[10][3] ), .B(\regZ[10][2] ), .Y(n4518) );
  NOR2X1 U2000 ( .A(\regZ[10][7] ), .B(\regZ[10][6] ), .Y(n4516) );
  NOR2X1 U2001 ( .A(\regZ[10][5] ), .B(\regZ[10][4] ), .Y(n4515) );
  NAND3X1 U2002 ( .A(n4519), .B(n4520), .C(n4521), .Y(n4325) );
  NOR2X1 U2003 ( .A(\regZ[9][1] ), .B(n4522), .Y(n4521) );
  OR2X1 U2004 ( .A(\regZ[9][3] ), .B(\regZ[9][2] ), .Y(n4522) );
  NOR2X1 U2005 ( .A(\regZ[9][7] ), .B(\regZ[9][6] ), .Y(n4520) );
  NOR2X1 U2006 ( .A(\regZ[9][5] ), .B(\regZ[9][4] ), .Y(n4519) );
  NAND2X1 U2007 ( .A(n4523), .B(n4524), .Y(n4502) );
  AOI22X1 U2008 ( .A(n4525), .B(n3827), .C(n3838), .D(n4329), .Y(n4524) );
  NAND3X1 U2009 ( .A(n4526), .B(n4527), .C(n4528), .Y(n4329) );
  NOR2X1 U2010 ( .A(\regZ[15][1] ), .B(n4529), .Y(n4528) );
  OR2X1 U2011 ( .A(\regZ[15][3] ), .B(\regZ[15][2] ), .Y(n4529) );
  NOR2X1 U2012 ( .A(\regZ[15][7] ), .B(\regZ[15][6] ), .Y(n4527) );
  NOR2X1 U2013 ( .A(\regZ[15][5] ), .B(\regZ[15][4] ), .Y(n4526) );
  AND2X1 U2014 ( .A(n4335), .B(n3583), .Y(n4525) );
  NAND3X1 U2015 ( .A(n4530), .B(n4531), .C(n4532), .Y(n4335) );
  NOR2X1 U2016 ( .A(\regZ[8][1] ), .B(n4533), .Y(n4532) );
  OR2X1 U2017 ( .A(\regZ[8][3] ), .B(\regZ[8][2] ), .Y(n4533) );
  NOR2X1 U2018 ( .A(\regZ[8][7] ), .B(\regZ[8][6] ), .Y(n4531) );
  NOR2X1 U2019 ( .A(\regZ[8][5] ), .B(\regZ[8][4] ), .Y(n4530) );
  AOI22X1 U2020 ( .A(n3865), .B(n4314), .C(n4480), .D(n4327), .Y(n4523) );
  NAND3X1 U2021 ( .A(n4534), .B(n4535), .C(n4536), .Y(n4327) );
  NOR2X1 U2022 ( .A(\regZ[13][1] ), .B(n4537), .Y(n4536) );
  OR2X1 U2023 ( .A(\regZ[13][3] ), .B(\regZ[13][2] ), .Y(n4537) );
  NOR2X1 U2024 ( .A(\regZ[13][7] ), .B(\regZ[13][6] ), .Y(n4535) );
  NOR2X1 U2025 ( .A(\regZ[13][5] ), .B(\regZ[13][4] ), .Y(n4534) );
  NAND3X1 U2026 ( .A(n4538), .B(n4539), .C(n4540), .Y(n4314) );
  NOR2X1 U2027 ( .A(\regZ[14][1] ), .B(n4541), .Y(n4540) );
  OR2X1 U2028 ( .A(\regZ[14][3] ), .B(\regZ[14][2] ), .Y(n4541) );
  NOR2X1 U2029 ( .A(\regZ[14][7] ), .B(\regZ[14][6] ), .Y(n4539) );
  NOR2X1 U2030 ( .A(\regZ[14][5] ), .B(\regZ[14][4] ), .Y(n4538) );
  INVX1 U2031 ( .A(n4542), .Y(n4364) );
  NAND3X1 U2032 ( .A(n4543), .B(n4544), .C(n4545), .Y(n4542) );
  NOR2X1 U2033 ( .A(\regZ[2][1] ), .B(n4546), .Y(n4545) );
  OR2X1 U2034 ( .A(\regZ[2][3] ), .B(\regZ[2][2] ), .Y(n4546) );
  NOR2X1 U2035 ( .A(\regZ[2][7] ), .B(\regZ[2][6] ), .Y(n4544) );
  NOR2X1 U2036 ( .A(\regZ[2][5] ), .B(\regZ[2][4] ), .Y(n4543) );
  OAI21X1 U2037 ( .A(n4547), .B(n4548), .C(n4549), .Y(n4499) );
  OAI21X1 U2038 ( .A(n4550), .B(n4551), .C(n4441), .Y(n4549) );
  INVX1 U2039 ( .A(n4552), .Y(n4551) );
  AOI22X1 U2040 ( .A(n4376), .B(n3924), .C(n4365), .D(n3583), .Y(n4552) );
  NAND3X1 U2041 ( .A(n4553), .B(n4554), .C(n4555), .Y(n4365) );
  NOR2X1 U2042 ( .A(\regZ[0][1] ), .B(n4556), .Y(n4555) );
  OR2X1 U2043 ( .A(\regZ[0][3] ), .B(\regZ[0][2] ), .Y(n4556) );
  NOR2X1 U2044 ( .A(\regZ[0][7] ), .B(\regZ[0][6] ), .Y(n4554) );
  NOR2X1 U2045 ( .A(\regZ[0][5] ), .B(\regZ[0][4] ), .Y(n4553) );
  NAND3X1 U2046 ( .A(n4557), .B(n4558), .C(n4559), .Y(n4376) );
  NOR2X1 U2047 ( .A(\regZ[1][1] ), .B(n4560), .Y(n4559) );
  OR2X1 U2048 ( .A(\regZ[1][3] ), .B(\regZ[1][2] ), .Y(n4560) );
  NOR2X1 U2049 ( .A(\regZ[1][7] ), .B(\regZ[1][6] ), .Y(n4558) );
  NOR2X1 U2050 ( .A(\regZ[1][5] ), .B(\regZ[1][4] ), .Y(n4557) );
  OAI21X1 U2051 ( .A(n4374), .B(n3641), .C(n4561), .Y(n4550) );
  AOI22X1 U2052 ( .A(n3865), .B(n4562), .C(n3838), .D(n4377), .Y(n4561) );
  NAND3X1 U2053 ( .A(n4565), .B(n4566), .C(n4567), .Y(n4377) );
  NOR2X1 U2054 ( .A(\regZ[7][1] ), .B(n4568), .Y(n4567) );
  OR2X1 U2055 ( .A(\regZ[7][3] ), .B(\regZ[7][2] ), .Y(n4568) );
  NOR2X1 U2056 ( .A(\regZ[7][7] ), .B(\regZ[7][6] ), .Y(n4566) );
  NOR2X1 U2057 ( .A(\regZ[7][5] ), .B(\regZ[7][4] ), .Y(n4565) );
  NAND3X1 U2058 ( .A(n4569), .B(n4570), .C(n4571), .Y(n4562) );
  NOR2X1 U2059 ( .A(\regZ[6][1] ), .B(n4575), .Y(n4571) );
  OR2X1 U2060 ( .A(\regZ[6][3] ), .B(\regZ[6][2] ), .Y(n4575) );
  NOR2X1 U2061 ( .A(\regZ[6][7] ), .B(\regZ[6][6] ), .Y(n4570) );
  NOR2X1 U2062 ( .A(\regZ[6][5] ), .B(\regZ[6][4] ), .Y(n4569) );
  INVX1 U2063 ( .A(n4576), .Y(n4374) );
  NAND3X1 U2064 ( .A(n4577), .B(n4578), .C(n4579), .Y(n4576) );
  NOR2X1 U2065 ( .A(\regZ[3][1] ), .B(n4580), .Y(n4579) );
  OR2X1 U2066 ( .A(\regZ[3][3] ), .B(\regZ[3][2] ), .Y(n4580) );
  NOR2X1 U2067 ( .A(\regZ[3][7] ), .B(\regZ[3][6] ), .Y(n4578) );
  NOR2X1 U2068 ( .A(\regZ[3][5] ), .B(\regZ[3][4] ), .Y(n4577) );
  NAND3X1 U2069 ( .A(n4581), .B(n4582), .C(n4583), .Y(n4548) );
  AOI22X1 U2070 ( .A(\regZ[2][0] ), .B(n4584), .C(\regZ[5][0] ), .D(n3877), 
        .Y(n4583) );
  INVX1 U2071 ( .A(n4438), .Y(n3877) );
  NAND2X1 U2072 ( .A(n4441), .B(n4480), .Y(n4438) );
  INVX1 U2073 ( .A(n3913), .Y(n4584) );
  NAND2X1 U2074 ( .A(n4441), .B(n4514), .Y(n3913) );
  NAND3X1 U2075 ( .A(n4441), .B(n3889), .C(\regZ[4][0] ), .Y(n4582) );
  OAI21X1 U2076 ( .A(n4585), .B(n4586), .C(n3586), .Y(n4581) );
  OAI21X1 U2077 ( .A(n3662), .B(n4587), .C(n4588), .Y(n4586) );
  AOI22X1 U2078 ( .A(\regZ[20][0] ), .B(n3889), .C(\regZ[19][0] ), .D(n3901), 
        .Y(n4588) );
  INVX1 U2079 ( .A(n3641), .Y(n3901) );
  INVX1 U2080 ( .A(\regZ[17][0] ), .Y(n4587) );
  NAND2X1 U2081 ( .A(n4589), .B(n4590), .Y(n4585) );
  AOI22X1 U2082 ( .A(n4591), .B(\regZ[16][0] ), .C(\regZ[23][0] ), .D(n3838), 
        .Y(n4590) );
  NOR2X1 U2083 ( .A(n3677), .B(n3585), .Y(n4591) );
  AOI22X1 U2084 ( .A(\regZ[22][0] ), .B(n3865), .C(\regZ[21][0] ), .D(n4480), 
        .Y(n4589) );
  NAND3X1 U2085 ( .A(n4592), .B(n4593), .C(n4594), .Y(n4547) );
  AOI22X1 U2086 ( .A(n4595), .B(\regZ[3][0] ), .C(n3585), .D(n4596), .Y(n4594)
         );
  NAND3X1 U2087 ( .A(n4597), .B(n4598), .C(n4599), .Y(n4596) );
  NOR2X1 U2088 ( .A(n4600), .B(n4601), .Y(n4599) );
  OAI21X1 U2089 ( .A(n3652), .B(n4602), .C(n4603), .Y(n4601) );
  MUX2X1 U2090 ( .B(n4604), .A(\regZ[24][0] ), .S(n3586), .Y(n4603) );
  NOR2X1 U2091 ( .A(n3677), .B(n4403), .Y(n4604) );
  INVX1 U2092 ( .A(\regZ[8][0] ), .Y(n4403) );
  INVX1 U2093 ( .A(\regZ[10][0] ), .Y(n4602) );
  OAI22X1 U2094 ( .A(n3662), .B(n4400), .C(n3641), .D(n4399), .Y(n4600) );
  INVX1 U2095 ( .A(\regZ[11][0] ), .Y(n4399) );
  INVX1 U2096 ( .A(\regZ[9][0] ), .Y(n4400) );
  AOI22X1 U2097 ( .A(\regZ[15][0] ), .B(n3838), .C(\regZ[14][0] ), .D(n3865), 
        .Y(n4598) );
  INVX1 U2098 ( .A(n3597), .Y(n3838) );
  AOI22X1 U2099 ( .A(\regZ[13][0] ), .B(n4480), .C(\regZ[12][0] ), .D(n3889), 
        .Y(n4597) );
  INVX1 U2100 ( .A(n3631), .Y(n3889) );
  NAND3X1 U2101 ( .A(n4605), .B(n4606), .C(n4607), .Y(n3631) );
  INVX1 U2102 ( .A(n3620), .Y(n4480) );
  NAND3X1 U2103 ( .A(n4606), .B(n4608), .C(n4605), .Y(n3620) );
  INVX1 U2104 ( .A(n3678), .Y(n3585) );
  NOR2X1 U2105 ( .A(n3641), .B(n3862), .Y(n4595) );
  NAND3X1 U2106 ( .A(n4609), .B(n4608), .C(n4610), .Y(n3641) );
  NAND3X1 U2107 ( .A(n4514), .B(n3586), .C(\regZ[18][0] ), .Y(n4593) );
  INVX1 U2108 ( .A(n3827), .Y(n3586) );
  INVX1 U2109 ( .A(n3652), .Y(n4514) );
  NAND3X1 U2110 ( .A(n4610), .B(n4609), .C(n4607), .Y(n3652) );
  OAI21X1 U2111 ( .A(n4611), .B(n4613), .C(n4441), .Y(n4592) );
  INVX1 U2112 ( .A(n3862), .Y(n4441) );
  NAND2X1 U2113 ( .A(n3827), .B(n3678), .Y(n3862) );
  XOR2X1 U2114 ( .A(n4614), .B(n4615), .Y(n3678) );
  XNOR2X1 U2115 ( .A(n4616), .B(n4617), .Y(n4614) );
  XOR2X1 U2116 ( .A(n4618), .B(n4619), .Y(n3827) );
  XNOR2X1 U2117 ( .A(n3940), .B(n3938), .Y(n4618) );
  AOI21X1 U2118 ( .A(n4616), .B(n4615), .C(n4628), .Y(n3938) );
  INVX1 U2119 ( .A(n4629), .Y(n4628) );
  OAI21X1 U2120 ( .A(n4615), .B(n4616), .C(n4617), .Y(n4629) );
  OAI21X1 U2121 ( .A(n4630), .B(n4631), .C(n4632), .Y(n4617) );
  OAI21X1 U2122 ( .A(n4633), .B(n4634), .C(n4635), .Y(n4632) );
  INVX1 U2123 ( .A(n4633), .Y(n4631) );
  AOI21X1 U2124 ( .A(n7204), .B(N3192), .C(n4682), .Y(n4615) );
  OAI21X1 U2125 ( .A(n4417), .B(n3943), .C(n4683), .Y(n4616) );
  INVX1 U2126 ( .A(n4421), .Y(n4417) );
  XOR2X1 U2127 ( .A(n4416), .B(n4415), .Y(n4421) );
  INVX1 U2128 ( .A(n4684), .Y(n4415) );
  XNOR2X1 U2129 ( .A(n4685), .B(n7204), .Y(n4416) );
  AOI21X1 U2130 ( .A(n7204), .B(N3193), .C(n4682), .Y(n3940) );
  INVX1 U2131 ( .A(n4686), .Y(n4613) );
  AOI22X1 U2132 ( .A(n3924), .B(\regZ[1][0] ), .C(n3583), .D(\regZ[0][0] ), 
        .Y(n4686) );
  INVX1 U2133 ( .A(n3677), .Y(n3583) );
  NAND3X1 U2134 ( .A(n4610), .B(n4605), .C(n4607), .Y(n3677) );
  INVX1 U2135 ( .A(n3662), .Y(n3924) );
  NAND3X1 U2136 ( .A(n4605), .B(n4608), .C(n4610), .Y(n3662) );
  OAI21X1 U2137 ( .A(n3597), .B(n4687), .C(n4688), .Y(n4611) );
  NAND2X1 U2138 ( .A(\regZ[6][0] ), .B(n3865), .Y(n4688) );
  INVX1 U2139 ( .A(n3609), .Y(n3865) );
  NAND3X1 U2140 ( .A(n4609), .B(n4606), .C(n4607), .Y(n3609) );
  INVX1 U2141 ( .A(\regZ[7][0] ), .Y(n4687) );
  NAND3X1 U2142 ( .A(n4606), .B(n4608), .C(n4609), .Y(n3597) );
  INVX1 U2143 ( .A(n4605), .Y(n4609) );
  XOR2X1 U2144 ( .A(n5089), .B(n5153), .Y(n4605) );
  XOR2X1 U2145 ( .A(n5154), .B(n5155), .Y(n5089) );
  INVX1 U2146 ( .A(n4607), .Y(n4608) );
  AOI21X1 U2147 ( .A(n5156), .B(n4408), .C(n5153), .Y(n4607) );
  INVX1 U2148 ( .A(n4610), .Y(n4606) );
  XOR2X1 U2149 ( .A(n5157), .B(n4633), .Y(n4610) );
  AOI21X1 U2150 ( .A(n7204), .B(N3191), .C(n4682), .Y(n4633) );
  XOR2X1 U2151 ( .A(n4635), .B(n4630), .Y(n5157) );
  INVX1 U2152 ( .A(n4634), .Y(n4630) );
  OAI21X1 U2153 ( .A(n5153), .B(n5158), .C(n5159), .Y(n4634) );
  OAI21X1 U2154 ( .A(n5154), .B(n5160), .C(n5155), .Y(n5159) );
  OAI21X1 U2155 ( .A(n5161), .B(n5162), .C(n5163), .Y(n5155) );
  AOI21X1 U2156 ( .A(n7204), .B(n4433), .C(n5164), .Y(n5163) );
  INVX1 U2157 ( .A(n5165), .Y(n5162) );
  INVX1 U2158 ( .A(n5153), .Y(n5160) );
  INVX1 U2159 ( .A(n5154), .Y(n5158) );
  AOI21X1 U2160 ( .A(n7204), .B(N3190), .C(n4682), .Y(n5154) );
  NOR2X1 U2161 ( .A(n4242), .B(n5161), .Y(n4682) );
  INVX1 U2162 ( .A(dx[1]), .Y(n4242) );
  NOR2X1 U2163 ( .A(n4408), .B(n5156), .Y(n5153) );
  AOI22X1 U2164 ( .A(dx[0]), .B(n7202), .C(n7204), .D(N3189), .Y(n5156) );
  INVX1 U2165 ( .A(n5166), .Y(n4408) );
  OAI21X1 U2166 ( .A(n7204), .B(n5167), .C(n5168), .Y(n5166) );
  INVX1 U2167 ( .A(n5169), .Y(n4635) );
  AOI22X1 U2168 ( .A(n5170), .B(n7202), .C(n4424), .D(n7204), .Y(n5169) );
  OAI21X1 U2169 ( .A(n4433), .B(n5171), .C(n4684), .Y(n4424) );
  NAND2X1 U2170 ( .A(n5171), .B(n4433), .Y(n4684) );
  XOR2X1 U2171 ( .A(n5172), .B(n3943), .Y(n5171) );
  INVX1 U2172 ( .A(n4436), .Y(n4433) );
  NAND2X1 U2173 ( .A(n5173), .B(n5168), .Y(n4436) );
  NAND2X1 U2174 ( .A(n5167), .B(n7204), .Y(n5168) );
  XOR2X1 U2175 ( .A(n7204), .B(n5174), .Y(n5167) );
  XOR2X1 U2176 ( .A(n3943), .B(n5175), .Y(n5173) );
  INVX1 U2177 ( .A(\Out_bThres[0] ), .Y(n4294) );
  MUX2X1 U2178 ( .B(n7716), .A(n5176), .S(n5177), .Y(n4651) );
  INVX1 U2179 ( .A(N4441), .Y(n7716) );
  OAI21X1 U2180 ( .A(n7717), .B(n5177), .C(n5178), .Y(n4650) );
  INVX1 U2181 ( .A(N4442), .Y(n7717) );
  OAI21X1 U2182 ( .A(n7718), .B(n5177), .C(n5179), .Y(n4649) );
  AND2X1 U2183 ( .A(n5180), .B(n5181), .Y(n5179) );
  INVX1 U2184 ( .A(N4438), .Y(n7718) );
  OAI21X1 U2185 ( .A(n7719), .B(n5177), .C(n5178), .Y(n4648) );
  INVX1 U2186 ( .A(N4439), .Y(n7719) );
  MUX2X1 U2187 ( .B(n7715), .A(n5176), .S(n5177), .Y(n4647) );
  INVX1 U2188 ( .A(N4435), .Y(n7715) );
  OAI21X1 U2189 ( .A(n7720), .B(n5177), .C(n5178), .Y(n4646) );
  INVX1 U2190 ( .A(N4436), .Y(n7720) );
  NAND2X1 U2191 ( .A(n5182), .B(n5181), .Y(n4645) );
  INVX1 U2192 ( .A(n5183), .Y(n5182) );
  MUX2X1 U2193 ( .B(n7721), .A(n5184), .S(n5177), .Y(n5183) );
  INVX1 U2194 ( .A(N4432), .Y(n7721) );
  OAI21X1 U2195 ( .A(n7722), .B(n5177), .C(n5178), .Y(n4644) );
  INVX1 U2196 ( .A(N4433), .Y(n7722) );
  OAI21X1 U2197 ( .A(n7723), .B(n5177), .C(n5181), .Y(n4643) );
  INVX1 U2198 ( .A(N4429), .Y(n7723) );
  OAI21X1 U2199 ( .A(n7724), .B(n5177), .C(n5178), .Y(n4642) );
  INVX1 U2200 ( .A(N4430), .Y(n7724) );
  MUX2X1 U2201 ( .B(n7725), .A(n5184), .S(n5177), .Y(n4641) );
  INVX1 U2202 ( .A(N4426), .Y(n7725) );
  OAI21X1 U2203 ( .A(n7726), .B(n5177), .C(n5178), .Y(n4640) );
  INVX1 U2204 ( .A(N4427), .Y(n7726) );
  OAI21X1 U2205 ( .A(n7727), .B(n5177), .C(n5181), .Y(n4639) );
  OAI21X1 U2206 ( .A(n5444), .B(n5445), .C(n5177), .Y(n5181) );
  NOR2X1 U2207 ( .A(n5446), .B(n5447), .Y(n5445) );
  OR2X1 U2208 ( .A(n5448), .B(\U3/U136/Z_0 ), .Y(n5447) );
  INVX1 U2209 ( .A(n5449), .Y(n5444) );
  INVX1 U2210 ( .A(N4423), .Y(n7727) );
  OAI21X1 U2211 ( .A(n7728), .B(n5177), .C(n5178), .Y(n4638) );
  INVX1 U2212 ( .A(N4424), .Y(n7728) );
  OAI21X1 U2213 ( .A(n7714), .B(n5177), .C(n5180), .Y(n4637) );
  OR2X1 U2214 ( .A(n5450), .B(n5451), .Y(n5180) );
  INVX1 U2215 ( .A(N4420), .Y(n7714) );
  OAI21X1 U2216 ( .A(n7729), .B(n5177), .C(n5178), .Y(n4636) );
  NAND2X1 U2217 ( .A(n5177), .B(n3557), .Y(n5178) );
  INVX1 U2218 ( .A(n5451), .Y(n5177) );
  NAND3X1 U2219 ( .A(n4131), .B(n5452), .C(n3936), .Y(n5451) );
  NAND3X1 U2220 ( .A(n5453), .B(n3548), .C(n5454), .Y(n5452) );
  OAI21X1 U2221 ( .A(n5455), .B(n5456), .C(n5457), .Y(n5454) );
  OAI21X1 U2222 ( .A(\U3/U136/Z_0 ), .B(n5446), .C(n5176), .Y(n5456) );
  AND2X1 U2223 ( .A(n5450), .B(n5184), .Y(n5176) );
  NAND3X1 U2224 ( .A(N2880), .B(n3864), .C(n4080), .Y(n5184) );
  NAND3X1 U2225 ( .A(N3336), .B(n4301), .C(N2841), .Y(n5450) );
  INVX1 U2226 ( .A(n5458), .Y(n4301) );
  INVX1 U2227 ( .A(N2945), .Y(n5446) );
  NAND2X1 U2228 ( .A(n5459), .B(n5449), .Y(n5455) );
  NAND2X1 U2229 ( .A(n5460), .B(N2874), .Y(n5449) );
  AOI21X1 U2230 ( .A(N2841), .B(N3336), .C(n5458), .Y(n5460) );
  OAI21X1 U2231 ( .A(n5448), .B(n4128), .C(n5458), .Y(n5459) );
  NAND2X1 U2232 ( .A(n4128), .B(n5461), .Y(n5458) );
  INVX1 U2233 ( .A(N2880), .Y(n5448) );
  INVX1 U2234 ( .A(N4421), .Y(n7729) );
  MUX2X1 U2235 ( .B(n7737), .A(n5462), .S(n3535), .Y(n4627) );
  AND2X1 U2236 ( .A(n5463), .B(n5464), .Y(n5462) );
  AOI21X1 U2237 ( .A(Out_direction[0]), .B(n5465), .C(n5466), .Y(n5464) );
  OAI21X1 U2238 ( .A(n5467), .B(n5468), .C(n5469), .Y(n5466) );
  NAND3X1 U2239 ( .A(n5470), .B(\Out_bThres[0] ), .C(dReadReg[2]), .Y(n5469)
         );
  INVX1 U2240 ( .A(n3537), .Y(n5470) );
  NAND3X1 U2241 ( .A(n5471), .B(n5472), .C(n5473), .Y(n3537) );
  INVX1 U2242 ( .A(dReadReg[3]), .Y(n5472) );
  NAND2X1 U2243 ( .A(dReadReg[1]), .B(dReadReg[0]), .Y(n5468) );
  OAI21X1 U2244 ( .A(n5474), .B(n5475), .C(n3539), .Y(n5467) );
  NAND2X1 U2245 ( .A(n5476), .B(n5477), .Y(n5475) );
  NOR2X1 U2246 ( .A(n5478), .B(n5479), .Y(n5477) );
  OAI21X1 U2247 ( .A(n3786), .B(n5480), .C(n5481), .Y(n5479) );
  AOI22X1 U2248 ( .A(n5482), .B(\regX[13][0] ), .C(n5483), .D(N1615), .Y(n5481) );
  INVX1 U2249 ( .A(n5484), .Y(n5482) );
  OAI21X1 U2250 ( .A(n5485), .B(n3653), .C(n5486), .Y(n5478) );
  AOI22X1 U2251 ( .A(n5487), .B(N1735), .C(n5488), .D(N1677), .Y(n5486) );
  INVX1 U2252 ( .A(n5489), .Y(n5487) );
  NOR2X1 U2253 ( .A(n5490), .B(n5491), .Y(n5476) );
  OAI21X1 U2254 ( .A(n3600), .B(n5492), .C(n5493), .Y(n5491) );
  AOI22X1 U2255 ( .A(n5494), .B(\regX[23][0] ), .C(n5495), .D(\regX[19][0] ), 
        .Y(n5493) );
  INVX1 U2256 ( .A(n5496), .Y(n5494) );
  OAI21X1 U2257 ( .A(n5497), .B(n3805), .C(n5498), .Y(n5490) );
  AOI22X1 U2258 ( .A(n5499), .B(\regX[15][0] ), .C(n5500), .D(\regX[21][0] ), 
        .Y(n5498) );
  INVX1 U2259 ( .A(n5501), .Y(n5499) );
  NAND3X1 U2260 ( .A(n5502), .B(n5503), .C(n5504), .Y(n5474) );
  NOR2X1 U2261 ( .A(n5505), .B(n5506), .Y(n5504) );
  OAI21X1 U2262 ( .A(n3860), .B(n3841), .C(n5507), .Y(n5506) );
  AOI22X1 U2263 ( .A(\regX[24][0] ), .B(n3582), .C(n5508), .D(\regX[20][0] ), 
        .Y(n5507) );
  OAI21X1 U2264 ( .A(n3840), .B(n3828), .C(n5509), .Y(n5505) );
  AOI22X1 U2265 ( .A(n5510), .B(\regX[18][0] ), .C(\regX[5][0] ), .D(n3876), 
        .Y(n5509) );
  NOR2X1 U2266 ( .A(n5511), .B(n5512), .Y(n5503) );
  OAI22X1 U2267 ( .A(n3676), .B(n3666), .C(n3890), .D(n3879), .Y(n5512) );
  OAI22X1 U2268 ( .A(n3902), .B(n3891), .C(n3941), .D(n3933), .Y(n5511) );
  AOI21X1 U2269 ( .A(\regX[8][0] ), .B(n5513), .C(n5514), .Y(n5502) );
  OAI22X1 U2270 ( .A(n3912), .B(n3903), .C(n3925), .D(n3914), .Y(n5514) );
  AOI22X1 U2271 ( .A(Out_gradient[0]), .B(n5515), .C(Out_gf[0]), .D(n5516), 
        .Y(n5463) );
  INVX1 U2272 ( .A(n5517), .Y(n5516) );
  INVX1 U2273 ( .A(N4489), .Y(n7737) );
  OAI21X1 U2274 ( .A(n5518), .B(n5519), .C(n5520), .Y(n4626) );
  MUX2X1 U2275 ( .B(N4486), .A(n5521), .S(n3535), .Y(n5520) );
  OAI21X1 U2276 ( .A(n5517), .B(n5522), .C(n5523), .Y(n5521) );
  AOI22X1 U2277 ( .A(Out_direction[1]), .B(n5465), .C(Out_gradient[1]), .D(
        n5515), .Y(n5523) );
  NOR2X1 U2278 ( .A(n5524), .B(n5525), .Y(n5518) );
  NAND2X1 U2279 ( .A(n5526), .B(n5527), .Y(n5525) );
  NOR2X1 U2280 ( .A(n5528), .B(n5529), .Y(n5527) );
  OAI21X1 U2281 ( .A(n3770), .B(n5484), .C(n5530), .Y(n5529) );
  AOI22X1 U2282 ( .A(n5500), .B(\regX[21][1] ), .C(\regX[9][1] ), .D(n3816), 
        .Y(n5530) );
  OAI21X1 U2283 ( .A(n3681), .B(n5501), .C(n5531), .Y(n5528) );
  AOI22X1 U2284 ( .A(n5495), .B(\regX[19][1] ), .C(n5532), .D(\regX[22][1] ), 
        .Y(n5531) );
  NOR2X1 U2285 ( .A(n5533), .B(n5534), .Y(n5526) );
  OAI21X1 U2286 ( .A(n3860), .B(n3843), .C(n5535), .Y(n5534) );
  AOI22X1 U2287 ( .A(n5488), .B(N1678), .C(\regX[17][1] ), .D(n3665), .Y(n5535) );
  OAI21X1 U2288 ( .A(n3758), .B(n5489), .C(n5536), .Y(n5533) );
  AOI22X1 U2289 ( .A(n5483), .B(N1616), .C(n5537), .D(\regX[11][1] ), .Y(n5536) );
  NAND3X1 U2290 ( .A(n5538), .B(n5539), .C(n5540), .Y(n5524) );
  NOR2X1 U2291 ( .A(n5541), .B(n5542), .Y(n5540) );
  OAI21X1 U2292 ( .A(n3589), .B(n5496), .C(n5543), .Y(n5542) );
  AOI22X1 U2293 ( .A(\regX[24][1] ), .B(n3582), .C(n5508), .D(\regX[20][1] ), 
        .Y(n5543) );
  OAI21X1 U2294 ( .A(n3840), .B(n3830), .C(n5544), .Y(n5541) );
  AOI22X1 U2295 ( .A(n5510), .B(\regX[18][1] ), .C(\regX[5][1] ), .D(n3876), 
        .Y(n5544) );
  NOR2X1 U2296 ( .A(n5545), .B(n5546), .Y(n5539) );
  OAI22X1 U2297 ( .A(n3676), .B(n3668), .C(n3890), .D(n3881), .Y(n5546) );
  OAI22X1 U2298 ( .A(n3902), .B(n3893), .C(n3941), .D(n3934), .Y(n5545) );
  AOI21X1 U2299 ( .A(\regX[8][1] ), .B(n5513), .C(n5547), .Y(n5538) );
  OAI22X1 U2300 ( .A(n3912), .B(n3905), .C(n3925), .D(n3916), .Y(n5547) );
  OAI21X1 U2301 ( .A(n5548), .B(n5519), .C(n5549), .Y(n4625) );
  MUX2X1 U2302 ( .B(N4483), .A(n5550), .S(n3535), .Y(n5549) );
  OAI21X1 U2303 ( .A(n5517), .B(n5551), .C(n5552), .Y(n5550) );
  AOI22X1 U2304 ( .A(Out_direction[2]), .B(n5465), .C(Out_gradient[2]), .D(
        n5515), .Y(n5552) );
  NOR2X1 U2305 ( .A(n5553), .B(n5554), .Y(n5548) );
  NAND2X1 U2306 ( .A(n5555), .B(n5556), .Y(n5554) );
  NOR2X1 U2307 ( .A(n5557), .B(n5558), .Y(n5556) );
  OAI21X1 U2308 ( .A(n3771), .B(n5484), .C(n5559), .Y(n5558) );
  AOI22X1 U2309 ( .A(n5500), .B(\regX[21][2] ), .C(\regX[9][2] ), .D(n3816), 
        .Y(n5559) );
  OAI21X1 U2310 ( .A(n3740), .B(n5501), .C(n5560), .Y(n5557) );
  AOI22X1 U2311 ( .A(n5495), .B(\regX[19][2] ), .C(n5532), .D(\regX[22][2] ), 
        .Y(n5560) );
  NOR2X1 U2312 ( .A(n5561), .B(n5562), .Y(n5555) );
  OAI21X1 U2313 ( .A(n3860), .B(n3844), .C(n5563), .Y(n5562) );
  AOI22X1 U2314 ( .A(n5488), .B(N1679), .C(\regX[17][2] ), .D(n3665), .Y(n5563) );
  OAI21X1 U2315 ( .A(n3759), .B(n5489), .C(n5564), .Y(n5561) );
  AOI22X1 U2316 ( .A(n5483), .B(N1617), .C(n5537), .D(\regX[11][2] ), .Y(n5564) );
  NAND3X1 U2317 ( .A(n5565), .B(n5566), .C(n5567), .Y(n5553) );
  NOR2X1 U2318 ( .A(n5568), .B(n5569), .Y(n5567) );
  OAI21X1 U2319 ( .A(n3590), .B(n5496), .C(n5570), .Y(n5569) );
  AOI22X1 U2320 ( .A(\regX[24][2] ), .B(n3582), .C(n5508), .D(\regX[20][2] ), 
        .Y(n5570) );
  OAI21X1 U2321 ( .A(n3840), .B(n3831), .C(n5571), .Y(n5568) );
  AOI22X1 U2322 ( .A(n5510), .B(\regX[18][2] ), .C(\regX[5][2] ), .D(n3876), 
        .Y(n5571) );
  NOR2X1 U2323 ( .A(n5572), .B(n5573), .Y(n5566) );
  OAI22X1 U2324 ( .A(n3676), .B(n3669), .C(n3890), .D(n3882), .Y(n5573) );
  OAI22X1 U2325 ( .A(n3902), .B(n3894), .C(n3941), .D(n3926), .Y(n5572) );
  AOI21X1 U2326 ( .A(\regX[8][2] ), .B(n5513), .C(n5574), .Y(n5565) );
  OAI22X1 U2327 ( .A(n3912), .B(n3906), .C(n3925), .D(n3917), .Y(n5574) );
  OAI21X1 U2328 ( .A(n5575), .B(n5519), .C(n5576), .Y(n4624) );
  MUX2X1 U2329 ( .B(N4480), .A(n5577), .S(n3535), .Y(n5576) );
  OAI21X1 U2330 ( .A(n5517), .B(n5578), .C(n5579), .Y(n5577) );
  AOI22X1 U2331 ( .A(Out_direction[3]), .B(n5465), .C(Out_gradient[3]), .D(
        n5515), .Y(n5579) );
  NOR2X1 U2332 ( .A(n5580), .B(n5581), .Y(n5575) );
  NAND2X1 U2333 ( .A(n5582), .B(n5583), .Y(n5581) );
  NOR2X1 U2334 ( .A(n5584), .B(n5585), .Y(n5583) );
  OAI21X1 U2335 ( .A(n3772), .B(n5484), .C(n5586), .Y(n5585) );
  AOI22X1 U2336 ( .A(n5500), .B(\regX[21][3] ), .C(\regX[9][3] ), .D(n3816), 
        .Y(n5586) );
  OAI21X1 U2337 ( .A(n3749), .B(n5501), .C(n5587), .Y(n5584) );
  AOI22X1 U2338 ( .A(n5495), .B(\regX[19][3] ), .C(n5532), .D(\regX[22][3] ), 
        .Y(n5587) );
  NOR2X1 U2339 ( .A(n5588), .B(n5589), .Y(n5582) );
  OAI21X1 U2340 ( .A(n3860), .B(n3845), .C(n5590), .Y(n5589) );
  AOI22X1 U2341 ( .A(n5488), .B(N1680), .C(\regX[17][3] ), .D(n3665), .Y(n5590) );
  OAI21X1 U2342 ( .A(n3760), .B(n5489), .C(n5591), .Y(n5588) );
  AOI22X1 U2343 ( .A(n5483), .B(N1618), .C(n5537), .D(\regX[11][3] ), .Y(n5591) );
  NAND3X1 U2344 ( .A(n5592), .B(n5593), .C(n5594), .Y(n5580) );
  NOR2X1 U2345 ( .A(n5595), .B(n5596), .Y(n5594) );
  OAI21X1 U2346 ( .A(n3591), .B(n5496), .C(n5597), .Y(n5596) );
  AOI22X1 U2347 ( .A(\regX[24][3] ), .B(n3582), .C(n5508), .D(\regX[20][3] ), 
        .Y(n5597) );
  OAI21X1 U2348 ( .A(n3840), .B(n3832), .C(n5598), .Y(n5595) );
  AOI22X1 U2349 ( .A(n5510), .B(\regX[18][3] ), .C(\regX[5][3] ), .D(n3876), 
        .Y(n5598) );
  NOR2X1 U2350 ( .A(n5599), .B(n5600), .Y(n5593) );
  OAI22X1 U2351 ( .A(n3676), .B(n3670), .C(n3890), .D(n3883), .Y(n5600) );
  OAI22X1 U2352 ( .A(n3902), .B(n3895), .C(n3941), .D(n3928), .Y(n5599) );
  AOI21X1 U2353 ( .A(\regX[8][3] ), .B(n5513), .C(n5601), .Y(n5592) );
  OAI22X1 U2354 ( .A(n3912), .B(n3907), .C(n3925), .D(n3918), .Y(n5601) );
  OAI21X1 U2355 ( .A(n5602), .B(n5519), .C(n5603), .Y(n4623) );
  MUX2X1 U2356 ( .B(N4477), .A(n5604), .S(n3535), .Y(n5603) );
  OAI21X1 U2357 ( .A(n5517), .B(n5605), .C(n5606), .Y(n5604) );
  AOI22X1 U2358 ( .A(Out_direction[4]), .B(n5465), .C(Out_gradient[4]), .D(
        n5515), .Y(n5606) );
  NOR2X1 U2359 ( .A(n5607), .B(n5608), .Y(n5602) );
  NAND2X1 U2360 ( .A(n5609), .B(n5610), .Y(n5608) );
  NOR2X1 U2361 ( .A(n5611), .B(n5612), .Y(n5610) );
  OAI21X1 U2362 ( .A(n3773), .B(n5484), .C(n5613), .Y(n5612) );
  AOI22X1 U2363 ( .A(n5500), .B(\regX[21][4] ), .C(\regX[9][4] ), .D(n3816), 
        .Y(n5613) );
  OAI21X1 U2364 ( .A(n3750), .B(n5501), .C(n5614), .Y(n5611) );
  AOI22X1 U2365 ( .A(n5495), .B(\regX[19][4] ), .C(n5532), .D(\regX[22][4] ), 
        .Y(n5614) );
  NOR2X1 U2366 ( .A(n5615), .B(n5616), .Y(n5609) );
  OAI21X1 U2367 ( .A(n3860), .B(n3846), .C(n5617), .Y(n5616) );
  AOI22X1 U2368 ( .A(n5488), .B(N1681), .C(\regX[17][4] ), .D(n3665), .Y(n5617) );
  OAI21X1 U2369 ( .A(n3761), .B(n5489), .C(n5618), .Y(n5615) );
  AOI22X1 U2370 ( .A(n5483), .B(N1619), .C(n5537), .D(\regX[11][4] ), .Y(n5618) );
  NAND3X1 U2371 ( .A(n5619), .B(n5620), .C(n5621), .Y(n5607) );
  NOR2X1 U2372 ( .A(n5622), .B(n5623), .Y(n5621) );
  OAI21X1 U2373 ( .A(n3592), .B(n5496), .C(n5624), .Y(n5623) );
  AOI22X1 U2374 ( .A(\regX[24][4] ), .B(n3582), .C(n5508), .D(\regX[20][4] ), 
        .Y(n5624) );
  OAI21X1 U2375 ( .A(n3840), .B(n3833), .C(n5625), .Y(n5622) );
  AOI22X1 U2376 ( .A(n5510), .B(\regX[18][4] ), .C(\regX[5][4] ), .D(n3876), 
        .Y(n5625) );
  NOR2X1 U2377 ( .A(n5626), .B(n5627), .Y(n5620) );
  OAI22X1 U2378 ( .A(n3676), .B(n3671), .C(n3890), .D(n3884), .Y(n5627) );
  INVX1 U2379 ( .A(\regX[16][4] ), .Y(n3671) );
  OAI22X1 U2380 ( .A(n3902), .B(n3896), .C(n3941), .D(n3929), .Y(n5626) );
  AOI21X1 U2381 ( .A(\regX[8][4] ), .B(n5513), .C(n5628), .Y(n5619) );
  OAI22X1 U2382 ( .A(n3912), .B(n3908), .C(n3925), .D(n3919), .Y(n5628) );
  OAI21X1 U2383 ( .A(n5629), .B(n5519), .C(n5630), .Y(n4622) );
  MUX2X1 U2384 ( .B(N4474), .A(n5631), .S(n3535), .Y(n5630) );
  OAI21X1 U2385 ( .A(n5517), .B(n5632), .C(n5633), .Y(n5631) );
  AOI22X1 U2386 ( .A(Out_direction[5]), .B(n5465), .C(Out_gradient[5]), .D(
        n5515), .Y(n5633) );
  NOR2X1 U2387 ( .A(n5634), .B(n5635), .Y(n5629) );
  NAND2X1 U2388 ( .A(n5636), .B(n5637), .Y(n5635) );
  NOR2X1 U2389 ( .A(n5638), .B(n5639), .Y(n5637) );
  OAI21X1 U2390 ( .A(n3774), .B(n5484), .C(n5640), .Y(n5639) );
  AOI22X1 U2391 ( .A(n5500), .B(\regX[21][5] ), .C(\regX[9][5] ), .D(n3816), 
        .Y(n5640) );
  OAI21X1 U2392 ( .A(n3751), .B(n5501), .C(n5641), .Y(n5638) );
  AOI22X1 U2393 ( .A(n5495), .B(\regX[19][5] ), .C(n5532), .D(\regX[22][5] ), 
        .Y(n5641) );
  NOR2X1 U2394 ( .A(n5642), .B(n5643), .Y(n5636) );
  OAI21X1 U2395 ( .A(n3860), .B(n3847), .C(n5644), .Y(n5643) );
  AOI22X1 U2396 ( .A(n5488), .B(N1682), .C(\regX[17][5] ), .D(n3665), .Y(n5644) );
  OAI21X1 U2397 ( .A(n3762), .B(n5489), .C(n5645), .Y(n5642) );
  AOI22X1 U2398 ( .A(n5483), .B(N1620), .C(n5537), .D(\regX[11][5] ), .Y(n5645) );
  NAND3X1 U2399 ( .A(n5646), .B(n5647), .C(n5648), .Y(n5634) );
  NOR2X1 U2400 ( .A(n5649), .B(n5650), .Y(n5648) );
  OAI21X1 U2401 ( .A(n3593), .B(n5496), .C(n5651), .Y(n5650) );
  AOI22X1 U2402 ( .A(\regX[24][5] ), .B(n3582), .C(n5508), .D(\regX[20][5] ), 
        .Y(n5651) );
  OAI21X1 U2403 ( .A(n3840), .B(n3834), .C(n5652), .Y(n5649) );
  AOI22X1 U2404 ( .A(n5510), .B(\regX[18][5] ), .C(\regX[5][5] ), .D(n3876), 
        .Y(n5652) );
  NOR2X1 U2405 ( .A(n5653), .B(n5654), .Y(n5647) );
  OAI22X1 U2406 ( .A(n3676), .B(n3672), .C(n3890), .D(n3885), .Y(n5654) );
  INVX1 U2407 ( .A(\regX[16][5] ), .Y(n3672) );
  OAI22X1 U2408 ( .A(n3902), .B(n3897), .C(n3941), .D(n3930), .Y(n5653) );
  AOI21X1 U2409 ( .A(\regX[8][5] ), .B(n5513), .C(n5655), .Y(n5646) );
  OAI22X1 U2410 ( .A(n3912), .B(n3909), .C(n3925), .D(n3920), .Y(n5655) );
  OAI21X1 U2411 ( .A(n5656), .B(n5519), .C(n5657), .Y(n4621) );
  MUX2X1 U2412 ( .B(N4471), .A(n5658), .S(n3535), .Y(n5657) );
  OAI21X1 U2413 ( .A(n5517), .B(n5659), .C(n5660), .Y(n5658) );
  AOI22X1 U2414 ( .A(Out_direction[6]), .B(n5465), .C(Out_gradient[6]), .D(
        n5515), .Y(n5660) );
  NOR2X1 U2415 ( .A(n5661), .B(n5662), .Y(n5656) );
  NAND2X1 U2416 ( .A(n5663), .B(n5664), .Y(n5662) );
  NOR2X1 U2417 ( .A(n5665), .B(n5666), .Y(n5664) );
  OAI21X1 U2418 ( .A(n3775), .B(n5484), .C(n5667), .Y(n5666) );
  AOI22X1 U2419 ( .A(n5500), .B(\regX[21][6] ), .C(\regX[9][6] ), .D(n3816), 
        .Y(n5667) );
  OAI21X1 U2420 ( .A(n3752), .B(n5501), .C(n5668), .Y(n5665) );
  AOI22X1 U2421 ( .A(n5495), .B(\regX[19][6] ), .C(n5532), .D(\regX[22][6] ), 
        .Y(n5668) );
  NOR2X1 U2422 ( .A(n5669), .B(n5670), .Y(n5663) );
  OAI21X1 U2423 ( .A(n3860), .B(n3848), .C(n5671), .Y(n5670) );
  AOI22X1 U2424 ( .A(n5488), .B(N1683), .C(\regX[17][6] ), .D(n3665), .Y(n5671) );
  OAI21X1 U2425 ( .A(n3763), .B(n5489), .C(n5672), .Y(n5669) );
  AOI22X1 U2426 ( .A(n5483), .B(N1621), .C(n5537), .D(\regX[11][6] ), .Y(n5672) );
  NAND3X1 U2427 ( .A(n5673), .B(n5674), .C(n5675), .Y(n5661) );
  NOR2X1 U2428 ( .A(n5676), .B(n5677), .Y(n5675) );
  OAI21X1 U2429 ( .A(n3594), .B(n5496), .C(n5678), .Y(n5677) );
  AOI22X1 U2430 ( .A(\regX[24][6] ), .B(n3582), .C(n5508), .D(\regX[20][6] ), 
        .Y(n5678) );
  OAI21X1 U2431 ( .A(n3840), .B(n3835), .C(n5679), .Y(n5676) );
  AOI22X1 U2432 ( .A(n5510), .B(\regX[18][6] ), .C(\regX[5][6] ), .D(n3876), 
        .Y(n5679) );
  NOR2X1 U2433 ( .A(n5680), .B(n5681), .Y(n5674) );
  OAI22X1 U2434 ( .A(n3676), .B(n3673), .C(n3890), .D(n3886), .Y(n5681) );
  INVX1 U2435 ( .A(\regX[16][6] ), .Y(n3673) );
  OAI22X1 U2436 ( .A(n3902), .B(n3898), .C(n3941), .D(n3931), .Y(n5680) );
  AOI21X1 U2437 ( .A(\regX[8][6] ), .B(n5513), .C(n5682), .Y(n5673) );
  OAI22X1 U2438 ( .A(n3912), .B(n3910), .C(n3925), .D(n3921), .Y(n5682) );
  OAI21X1 U2439 ( .A(n5683), .B(n5519), .C(n5684), .Y(n4620) );
  MUX2X1 U2440 ( .B(N4468), .A(n5685), .S(n3535), .Y(n5684) );
  OAI21X1 U2441 ( .A(n5517), .B(n5686), .C(n5687), .Y(n5685) );
  AOI22X1 U2442 ( .A(Out_direction[7]), .B(n5465), .C(Out_gradient[7]), .D(
        n5515), .Y(n5687) );
  INVX1 U2443 ( .A(n5688), .Y(n5515) );
  NAND3X1 U2444 ( .A(n3539), .B(n5471), .C(dReadReg[0]), .Y(n5688) );
  INVX1 U2445 ( .A(n5689), .Y(n5465) );
  NAND3X1 U2446 ( .A(n3539), .B(n5473), .C(dReadReg[1]), .Y(n5689) );
  NAND3X1 U2447 ( .A(n5473), .B(n5471), .C(n3539), .Y(n5517) );
  NAND3X1 U2448 ( .A(n3539), .B(n3535), .C(n5690), .Y(n5519) );
  NOR2X1 U2449 ( .A(n5473), .B(n5471), .Y(n5690) );
  INVX1 U2450 ( .A(dReadReg[1]), .Y(n5471) );
  INVX1 U2451 ( .A(dReadReg[0]), .Y(n5473) );
  INVX1 U2452 ( .A(n5691), .Y(n3535) );
  NAND3X1 U2453 ( .A(rst_b), .B(n5692), .C(bWE), .Y(n5691) );
  NOR2X1 U2454 ( .A(dReadReg[2]), .B(dReadReg[3]), .Y(n3539) );
  NOR2X1 U2455 ( .A(n5693), .B(n5694), .Y(n5683) );
  NAND2X1 U2456 ( .A(n5695), .B(n5696), .Y(n5694) );
  NOR2X1 U2457 ( .A(n5697), .B(n5698), .Y(n5696) );
  OAI21X1 U2458 ( .A(n3767), .B(n5484), .C(n5699), .Y(n5698) );
  AOI22X1 U2459 ( .A(n5500), .B(\regX[21][7] ), .C(\regX[9][7] ), .D(n3816), 
        .Y(n5699) );
  INVX1 U2460 ( .A(n5497), .Y(n3816) );
  NAND2X1 U2461 ( .A(n4195), .B(n5700), .Y(n5497) );
  AND2X1 U2462 ( .A(n3785), .B(n4181), .Y(n5500) );
  NAND2X1 U2463 ( .A(n4195), .B(n3785), .Y(n5484) );
  OAI21X1 U2464 ( .A(n3753), .B(n5501), .C(n5701), .Y(n5697) );
  AOI22X1 U2465 ( .A(n5495), .B(\regX[19][7] ), .C(n5532), .D(\regX[22][7] ), 
        .Y(n5701) );
  INVX1 U2466 ( .A(n5492), .Y(n5532) );
  NAND2X1 U2467 ( .A(n4183), .B(n3766), .Y(n5492) );
  AND2X1 U2468 ( .A(n3804), .B(n4181), .Y(n5495) );
  NAND2X1 U2469 ( .A(n4195), .B(n3766), .Y(n5501) );
  NOR2X1 U2470 ( .A(n5702), .B(n5703), .Y(n5695) );
  OAI21X1 U2471 ( .A(n3860), .B(n3849), .C(n5704), .Y(n5703) );
  AOI22X1 U2472 ( .A(n5488), .B(N1684), .C(\regX[17][7] ), .D(n3665), .Y(n5704) );
  INVX1 U2473 ( .A(n5485), .Y(n3665) );
  NAND2X1 U2474 ( .A(n4181), .B(n5700), .Y(n5485) );
  AND2X1 U2475 ( .A(n4197), .B(n3785), .Y(n5488) );
  OAI21X1 U2476 ( .A(n3764), .B(n5489), .C(n5705), .Y(n5702) );
  AOI22X1 U2477 ( .A(n5483), .B(N1622), .C(n5537), .D(\regX[11][7] ), .Y(n5705) );
  INVX1 U2478 ( .A(n5480), .Y(n5537) );
  NAND2X1 U2479 ( .A(n4195), .B(n3804), .Y(n5480) );
  NOR2X1 U2480 ( .A(n5706), .B(n3664), .Y(n4195) );
  AND2X1 U2481 ( .A(n4197), .B(n3804), .Y(n5483) );
  NAND2X1 U2482 ( .A(n4197), .B(n3766), .Y(n5489) );
  NOR2X1 U2483 ( .A(n3664), .B(N977), .Y(n4197) );
  NAND3X1 U2484 ( .A(n5707), .B(n5708), .C(n5709), .Y(n5693) );
  NOR2X1 U2485 ( .A(n5710), .B(n5711), .Y(n5709) );
  OAI21X1 U2486 ( .A(n3595), .B(n5496), .C(n5712), .Y(n5711) );
  AOI22X1 U2487 ( .A(\regX[24][7] ), .B(n3582), .C(n5508), .D(\regX[20][7] ), 
        .Y(n5712) );
  AND2X1 U2488 ( .A(n3785), .B(n4183), .Y(n5508) );
  NOR2X1 U2489 ( .A(n3815), .B(n3664), .Y(n3582) );
  NAND2X1 U2490 ( .A(n4181), .B(n3766), .Y(n5496) );
  NOR2X1 U2491 ( .A(n5706), .B(n3815), .Y(n4181) );
  OAI21X1 U2492 ( .A(n3840), .B(n3836), .C(n5713), .Y(n5710) );
  AOI22X1 U2493 ( .A(n5510), .B(\regX[18][7] ), .C(\regX[5][7] ), .D(n3876), 
        .Y(n5713) );
  INVX1 U2494 ( .A(n4204), .Y(n3876) );
  NAND2X1 U2495 ( .A(n5714), .B(n3785), .Y(n4204) );
  AND2X1 U2496 ( .A(n3804), .B(n4183), .Y(n5510) );
  NOR2X1 U2497 ( .A(n3815), .B(N977), .Y(n4183) );
  NAND2X1 U2498 ( .A(n5714), .B(n3766), .Y(n3840) );
  NOR2X1 U2499 ( .A(n5715), .B(n5716), .Y(n5708) );
  OAI22X1 U2500 ( .A(n3676), .B(n3674), .C(n3890), .D(n3887), .Y(n5716) );
  NAND2X1 U2501 ( .A(n3785), .B(n5717), .Y(n3890) );
  NOR2X1 U2502 ( .A(n5718), .B(N978), .Y(n3785) );
  INVX1 U2503 ( .A(\regX[16][7] ), .Y(n3674) );
  NAND3X1 U2504 ( .A(N981), .B(n3664), .C(n3580), .Y(n3676) );
  INVX1 U2505 ( .A(N980), .Y(n3664) );
  OAI22X1 U2506 ( .A(n3902), .B(n3899), .C(n3941), .D(n3932), .Y(n5715) );
  NAND2X1 U2507 ( .A(n3580), .B(n5719), .Y(n3941) );
  NAND2X1 U2508 ( .A(n5714), .B(n3804), .Y(n3902) );
  AOI21X1 U2509 ( .A(\regX[8][7] ), .B(n5513), .C(n5720), .Y(n5707) );
  OAI22X1 U2510 ( .A(n3912), .B(n3911), .C(n3925), .D(n3922), .Y(n5720) );
  NAND2X1 U2511 ( .A(n5714), .B(n5700), .Y(n3925) );
  AND2X1 U2512 ( .A(N977), .B(n5719), .Y(n5714) );
  NAND2X1 U2513 ( .A(n3804), .B(n5717), .Y(n3912) );
  NOR2X1 U2514 ( .A(n5721), .B(N979), .Y(n3804) );
  INVX1 U2515 ( .A(n3826), .Y(n5513) );
  NAND3X1 U2516 ( .A(N980), .B(n3815), .C(n3580), .Y(n3826) );
  AND2X1 U2517 ( .A(n5700), .B(n5706), .Y(n3580) );
  NOR2X1 U2518 ( .A(N979), .B(N978), .Y(n5700) );
  INVX1 U2519 ( .A(N981), .Y(n3815) );
  OR2X1 U2520 ( .A(bCE), .B(dAddrRegRow[0]), .Y(n4574) );
  OR2X1 U2521 ( .A(bCE), .B(dAddrRegRow[1]), .Y(n4573) );
  AND2X1 U2522 ( .A(dAddrRegRow[2]), .B(n5692), .Y(n4572) );
  MUX2X1 U2523 ( .B(n5722), .A(n4275), .S(n5723), .Y(n3748) );
  INVX1 U2524 ( .A(tpSum[7]), .Y(n4275) );
  INVX1 U2525 ( .A(Out_gf[0]), .Y(n5722) );
  MUX2X1 U2526 ( .B(n5522), .A(n4278), .S(n5723), .Y(n3747) );
  INVX1 U2527 ( .A(tpSum[8]), .Y(n4278) );
  INVX1 U2528 ( .A(Out_gf[1]), .Y(n5522) );
  MUX2X1 U2529 ( .B(n5551), .A(n4280), .S(n5723), .Y(n3746) );
  INVX1 U2530 ( .A(tpSum[9]), .Y(n4280) );
  INVX1 U2531 ( .A(Out_gf[2]), .Y(n5551) );
  MUX2X1 U2532 ( .B(n5578), .A(n4282), .S(n5723), .Y(n3745) );
  INVX1 U2533 ( .A(tpSum[10]), .Y(n4282) );
  INVX1 U2534 ( .A(Out_gf[3]), .Y(n5578) );
  MUX2X1 U2535 ( .B(n5605), .A(n4284), .S(n5723), .Y(n3744) );
  INVX1 U2536 ( .A(tpSum[11]), .Y(n4284) );
  INVX1 U2537 ( .A(Out_gf[4]), .Y(n5605) );
  MUX2X1 U2538 ( .B(n5632), .A(n4286), .S(n5723), .Y(n3743) );
  INVX1 U2539 ( .A(tpSum[12]), .Y(n4286) );
  INVX1 U2540 ( .A(Out_gf[5]), .Y(n5632) );
  MUX2X1 U2541 ( .B(n5659), .A(n4288), .S(n5723), .Y(n3742) );
  INVX1 U2542 ( .A(tpSum[13]), .Y(n4288) );
  INVX1 U2543 ( .A(Out_gf[6]), .Y(n5659) );
  MUX2X1 U2544 ( .B(n5686), .A(n4290), .S(n5723), .Y(n3741) );
  NOR2X1 U2545 ( .A(n4292), .B(n5453), .Y(n5723) );
  NAND3X1 U2546 ( .A(n3936), .B(n4250), .C(n5724), .Y(n4292) );
  INVX1 U2547 ( .A(n3850), .Y(n3936) );
  NAND2X1 U2548 ( .A(n3545), .B(rst_b), .Y(n3850) );
  INVX1 U2549 ( .A(tpSum[14]), .Y(n4290) );
  INVX1 U2550 ( .A(Out_gf[7]), .Y(n5686) );
  OAI22X1 U2551 ( .A(n3946), .B(n5726), .C(n3478), .D(n5727), .Y(n3739) );
  INVX1 U2552 ( .A(N2300), .Y(n5727) );
  OAI22X1 U2553 ( .A(n3946), .B(n5728), .C(n3478), .D(n5729), .Y(n3738) );
  INVX1 U2554 ( .A(N2301), .Y(n5729) );
  OAI22X1 U2555 ( .A(n3946), .B(n5730), .C(n3478), .D(n5731), .Y(n3737) );
  INVX1 U2556 ( .A(N2302), .Y(n5731) );
  OAI22X1 U2557 ( .A(n3946), .B(n5732), .C(n3478), .D(n5733), .Y(n3736) );
  INVX1 U2558 ( .A(N2303), .Y(n5733) );
  OAI22X1 U2559 ( .A(n3946), .B(n5734), .C(n3478), .D(n5735), .Y(n3735) );
  INVX1 U2560 ( .A(N2304), .Y(n5735) );
  OAI22X1 U2561 ( .A(n3946), .B(n5736), .C(n3478), .D(n5737), .Y(n3734) );
  INVX1 U2562 ( .A(N2305), .Y(n5737) );
  OAI22X1 U2563 ( .A(n3946), .B(n5738), .C(n4012), .D(n5739), .Y(n3733) );
  INVX1 U2564 ( .A(N2306), .Y(n5739) );
  OAI22X1 U2565 ( .A(n3946), .B(n5740), .C(n4012), .D(n5741), .Y(n3732) );
  INVX1 U2566 ( .A(N2307), .Y(n5741) );
  OAI22X1 U2567 ( .A(n3946), .B(n5742), .C(n4012), .D(n5743), .Y(n3731) );
  INVX1 U2568 ( .A(N2308), .Y(n5743) );
  OAI22X1 U2569 ( .A(n3946), .B(n5744), .C(n4012), .D(n5745), .Y(n3730) );
  INVX1 U2570 ( .A(N2309), .Y(n5745) );
  OAI22X1 U2571 ( .A(n3946), .B(n5746), .C(n4012), .D(n5747), .Y(n3729) );
  INVX1 U2572 ( .A(N2310), .Y(n5747) );
  OAI22X1 U2573 ( .A(n3946), .B(n5748), .C(n4012), .D(n5749), .Y(n3728) );
  INVX1 U2574 ( .A(N2311), .Y(n5749) );
  OAI22X1 U2575 ( .A(n3946), .B(n5750), .C(n4012), .D(n5751), .Y(n3727) );
  INVX1 U2576 ( .A(N2312), .Y(n5751) );
  OAI22X1 U2577 ( .A(n3946), .B(n5752), .C(n4012), .D(n5753), .Y(n3726) );
  INVX1 U2578 ( .A(N2313), .Y(n5753) );
  OAI22X1 U2579 ( .A(n3946), .B(n5754), .C(n4012), .D(n5755), .Y(n3725) );
  INVX1 U2580 ( .A(N2314), .Y(n5755) );
  OAI22X1 U2581 ( .A(n3946), .B(n5756), .C(n4012), .D(n5757), .Y(n3724) );
  INVX1 U2582 ( .A(N2315), .Y(n5757) );
  OAI22X1 U2583 ( .A(n3946), .B(n5758), .C(n4012), .D(n5759), .Y(n3723) );
  INVX1 U2584 ( .A(N2316), .Y(n5759) );
  OAI22X1 U2585 ( .A(n3946), .B(n5760), .C(n4012), .D(n5761), .Y(n3722) );
  INVX1 U2586 ( .A(N2317), .Y(n5761) );
  OAI22X1 U2587 ( .A(n3946), .B(n5762), .C(n4012), .D(n5763), .Y(n3721) );
  INVX1 U2588 ( .A(N2318), .Y(n5763) );
  OAI22X1 U2589 ( .A(n3946), .B(n5764), .C(n4012), .D(n5765), .Y(n3720) );
  INVX1 U2590 ( .A(N2319), .Y(n5765) );
  OAI22X1 U2591 ( .A(n3946), .B(n5766), .C(n4012), .D(n5767), .Y(n3719) );
  INVX1 U2592 ( .A(N2320), .Y(n5767) );
  OAI22X1 U2593 ( .A(n3946), .B(n5768), .C(n4012), .D(n5769), .Y(n3718) );
  INVX1 U2594 ( .A(N2321), .Y(n5769) );
  OAI22X1 U2595 ( .A(n3946), .B(n5770), .C(n4012), .D(n5771), .Y(n3717) );
  INVX1 U2596 ( .A(N2322), .Y(n5771) );
  OAI22X1 U2597 ( .A(n3946), .B(n5772), .C(n4012), .D(n5773), .Y(n3716) );
  INVX1 U2598 ( .A(N2323), .Y(n5773) );
  OAI22X1 U2599 ( .A(n3946), .B(n5774), .C(n4012), .D(n5775), .Y(n3715) );
  INVX1 U2600 ( .A(N2324), .Y(n5775) );
  OAI22X1 U2601 ( .A(n3946), .B(n5776), .C(n4012), .D(n5777), .Y(n3714) );
  INVX1 U2602 ( .A(N2325), .Y(n5777) );
  OAI22X1 U2603 ( .A(n3946), .B(n5778), .C(n4012), .D(n5779), .Y(n3713) );
  INVX1 U2604 ( .A(N2326), .Y(n5779) );
  OAI22X1 U2605 ( .A(n3946), .B(n5780), .C(n4012), .D(n5781), .Y(n3712) );
  INVX1 U2606 ( .A(N2327), .Y(n5781) );
  OAI22X1 U2607 ( .A(n3946), .B(n5782), .C(n4012), .D(n5783), .Y(n3711) );
  INVX1 U2608 ( .A(N2328), .Y(n5783) );
  OAI22X1 U2609 ( .A(n3946), .B(n5784), .C(n4012), .D(n5785), .Y(n3710) );
  INVX1 U2610 ( .A(N2329), .Y(n5785) );
  OAI22X1 U2611 ( .A(n3946), .B(n5786), .C(n4012), .D(n5787), .Y(n3709) );
  INVX1 U2612 ( .A(N2330), .Y(n5787) );
  OAI22X1 U2613 ( .A(n3946), .B(n5788), .C(n4012), .D(n5789), .Y(n3708) );
  INVX1 U2614 ( .A(N2331), .Y(n5789) );
  NAND3X1 U2615 ( .A(n4257), .B(rst_b), .C(n3557), .Y(n4012) );
  NAND3X1 U2616 ( .A(rst_b), .B(n5453), .C(n3557), .Y(n5790) );
  AND2X1 U2617 ( .A(n3545), .B(n4273), .Y(n3557) );
  NAND2X1 U2618 ( .A(n3481), .B(n3476), .Y(n4273) );
  NOR2X1 U2619 ( .A(n5692), .B(bOPEnable), .Y(n3545) );
  INVX1 U2620 ( .A(n5792), .Y(n3706) );
  MUX2X1 U2621 ( .B(Gx[0]), .A(N2558), .S(n4272), .Y(n5792) );
  INVX1 U2622 ( .A(n5793), .Y(n3705) );
  MUX2X1 U2623 ( .B(Gx[1]), .A(N2559), .S(n4272), .Y(n5793) );
  INVX1 U2624 ( .A(n5794), .Y(n3704) );
  MUX2X1 U2625 ( .B(Gx[2]), .A(N2560), .S(n4272), .Y(n5794) );
  INVX1 U2626 ( .A(n5795), .Y(n3703) );
  MUX2X1 U2627 ( .B(Gx[3]), .A(N2561), .S(n4272), .Y(n5795) );
  INVX1 U2628 ( .A(n5796), .Y(n3702) );
  MUX2X1 U2629 ( .B(Gx[4]), .A(N2562), .S(n4272), .Y(n5796) );
  INVX1 U2630 ( .A(n5797), .Y(n3701) );
  MUX2X1 U2631 ( .B(Gx[5]), .A(N2563), .S(n4272), .Y(n5797) );
  INVX1 U2632 ( .A(n5798), .Y(n3700) );
  MUX2X1 U2633 ( .B(Gx[6]), .A(N2564), .S(n4272), .Y(n5798) );
  INVX1 U2634 ( .A(n5799), .Y(n3699) );
  MUX2X1 U2635 ( .B(Gx[7]), .A(N2565), .S(n4272), .Y(n5799) );
  INVX1 U2636 ( .A(n5800), .Y(n3698) );
  MUX2X1 U2637 ( .B(Gx[8]), .A(N2566), .S(n4272), .Y(n5800) );
  INVX1 U2638 ( .A(n5801), .Y(n3697) );
  MUX2X1 U2639 ( .B(Gx[9]), .A(N2567), .S(n4272), .Y(n5801) );
  INVX1 U2640 ( .A(n5802), .Y(n3696) );
  MUX2X1 U2641 ( .B(Gx[10]), .A(N2568), .S(n4272), .Y(n5802) );
  INVX1 U2642 ( .A(n5803), .Y(n3695) );
  MUX2X1 U2643 ( .B(N971), .A(N3189), .S(bCE), .Y(n5803) );
  INVX1 U2644 ( .A(n5804), .Y(n3694) );
  MUX2X1 U2645 ( .B(N972), .A(N3190), .S(bCE), .Y(n5804) );
  INVX1 U2646 ( .A(n5805), .Y(n3693) );
  MUX2X1 U2647 ( .B(N973), .A(N3191), .S(bCE), .Y(n5805) );
  INVX1 U2648 ( .A(n5806), .Y(n3692) );
  MUX2X1 U2649 ( .B(N974), .A(N3192), .S(bCE), .Y(n5806) );
  INVX1 U2650 ( .A(n5807), .Y(n3691) );
  MUX2X1 U2651 ( .B(N975), .A(N3193), .S(bCE), .Y(n5807) );
  INVX1 U2652 ( .A(n5808), .Y(n3690) );
  MUX2X1 U2653 ( .B(dAddrRegCol[2]), .A(n5170), .S(bCE), .Y(n5808) );
  OAI21X1 U2654 ( .A(n5165), .B(n5809), .C(n5810), .Y(n5170) );
  MUX2X1 U2655 ( .B(n5811), .A(n5812), .S(bCE), .Y(n3689) );
  NOR2X1 U2656 ( .A(n5164), .B(n5165), .Y(n5812) );
  NOR2X1 U2657 ( .A(n5175), .B(n5174), .Y(n5164) );
  INVX1 U2658 ( .A(dAddrRegCol[1]), .Y(n5811) );
  MUX2X1 U2659 ( .B(n4240), .A(n5813), .S(n3486), .Y(n3688) );
  INVX1 U2660 ( .A(InData[7]), .Y(n5813) );
  INVX1 U2661 ( .A(\regY[6][7] ), .Y(n4240) );
  MUX2X1 U2662 ( .B(n4233), .A(n5814), .S(n3486), .Y(n3687) );
  INVX1 U2663 ( .A(InData[5]), .Y(n5814) );
  INVX1 U2664 ( .A(\regY[6][5] ), .Y(n4233) );
  MUX2X1 U2665 ( .B(n4248), .A(n5815), .S(n3486), .Y(n3686) );
  INVX1 U2666 ( .A(InData[4]), .Y(n5815) );
  INVX1 U2667 ( .A(\regY[6][4] ), .Y(n4248) );
  MUX2X1 U2668 ( .B(n4253), .A(n5816), .S(n3486), .Y(n3685) );
  INVX1 U2669 ( .A(InData[3]), .Y(n5816) );
  INVX1 U2670 ( .A(\regY[6][3] ), .Y(n4253) );
  MUX2X1 U2671 ( .B(n4239), .A(n5817), .S(n3486), .Y(n3684) );
  INVX1 U2672 ( .A(InData[2]), .Y(n5817) );
  INVX1 U2673 ( .A(\regY[6][2] ), .Y(n4239) );
  MUX2X1 U2674 ( .B(n4237), .A(n5818), .S(n3486), .Y(n3683) );
  INVX1 U2675 ( .A(InData[1]), .Y(n5818) );
  INVX1 U2676 ( .A(\regY[6][1] ), .Y(n4237) );
  MUX2X1 U2677 ( .B(n4241), .A(n5819), .S(n3486), .Y(n3682) );
  NOR2X1 U2678 ( .A(n5820), .B(n5821), .Y(n3486) );
  NAND3X1 U2679 ( .A(n3490), .B(n3853), .C(n5822), .Y(n5821) );
  AND2X1 U2680 ( .A(dWriteReg[0]), .B(rst_b), .Y(n5822) );
  NOR2X1 U2681 ( .A(N983), .B(N982), .Y(n3853) );
  NOR2X1 U2682 ( .A(bCE), .B(bWE), .Y(n3490) );
  NAND3X1 U2683 ( .A(n3854), .B(n3944), .C(n4214), .Y(n5820) );
  NOR2X1 U2684 ( .A(dWriteReg[3]), .B(dWriteReg[2]), .Y(n4214) );
  INVX1 U2685 ( .A(dWriteReg[1]), .Y(n3944) );
  INVX1 U2686 ( .A(n3860), .Y(n3854) );
  NAND2X1 U2687 ( .A(n3766), .B(n5717), .Y(n3860) );
  AND2X1 U2688 ( .A(n5719), .B(n5706), .Y(n5717) );
  INVX1 U2689 ( .A(N977), .Y(n5706) );
  NOR2X1 U2690 ( .A(N981), .B(N980), .Y(n5719) );
  NOR2X1 U2691 ( .A(n5718), .B(n5721), .Y(n3766) );
  INVX1 U2692 ( .A(N978), .Y(n5721) );
  INVX1 U2693 ( .A(N979), .Y(n5718) );
  INVX1 U2694 ( .A(InData[0]), .Y(n5819) );
  INVX1 U2695 ( .A(\regY[6][0] ), .Y(n4241) );
  NAND2X1 U2696 ( .A(n3475), .B(n3476), .Y(n2980) );
  OAI21X1 U2697 ( .A(n3475), .B(n3619), .C(n5824), .Y(\U3/U98/Z_7 ) );
  OAI21X1 U2698 ( .A(n3475), .B(n3618), .C(n5824), .Y(\U3/U98/Z_6 ) );
  OAI21X1 U2699 ( .A(n3475), .B(n3617), .C(n5824), .Y(\U3/U98/Z_5 ) );
  OAI21X1 U2700 ( .A(n3475), .B(n3616), .C(n5824), .Y(\U3/U98/Z_4 ) );
  OAI21X1 U2701 ( .A(n3475), .B(n3615), .C(n5824), .Y(\U3/U98/Z_3 ) );
  OAI21X1 U2702 ( .A(n3475), .B(n3614), .C(n5824), .Y(\U3/U98/Z_2 ) );
  OAI21X1 U2703 ( .A(n3475), .B(n3613), .C(n5824), .Y(\U3/U98/Z_1 ) );
  NAND2X1 U2704 ( .A(dy[1]), .B(n7204), .Y(n5824) );
  OAI22X1 U2705 ( .A(n3943), .B(n5825), .C(n3475), .D(n3611), .Y(\U3/U98/Z_0 )
         );
  NAND2X1 U2706 ( .A(n3943), .B(n3475), .Y(\U3/U97/Z_0 ) );
  NAND2X1 U2707 ( .A(n3481), .B(n3482), .Y(\U3/U96/Z_0 ) );
  NAND2X1 U2708 ( .A(n5827), .B(n3482), .Y(\U3/U95/Z_0 ) );
  AND2X1 U2709 ( .A(N2890), .B(n7240), .Y(\U3/U94/Z_9 ) );
  AND2X1 U2710 ( .A(N2889), .B(n7240), .Y(\U3/U94/Z_8 ) );
  OAI21X1 U2711 ( .A(n5827), .B(n3849), .C(n5828), .Y(\U3/U94/Z_7 ) );
  NAND2X1 U2712 ( .A(N2888), .B(n7240), .Y(n5828) );
  OAI21X1 U2713 ( .A(n5827), .B(n3848), .C(n5829), .Y(\U3/U94/Z_6 ) );
  NAND2X1 U2714 ( .A(N2887), .B(n7240), .Y(n5829) );
  OAI21X1 U2715 ( .A(n5827), .B(n3847), .C(n5830), .Y(\U3/U94/Z_5 ) );
  NAND2X1 U2716 ( .A(N2886), .B(n7240), .Y(n5830) );
  OAI21X1 U2717 ( .A(n5827), .B(n3846), .C(n5831), .Y(\U3/U94/Z_4 ) );
  NAND2X1 U2718 ( .A(N2885), .B(n7240), .Y(n5831) );
  NOR2X1 U2719 ( .A(n3482), .B(n5832), .Y(\U3/U94/Z_31 ) );
  OAI21X1 U2720 ( .A(n3845), .B(n5827), .C(n5833), .Y(\U3/U94/Z_3 ) );
  NAND2X1 U2721 ( .A(N2884), .B(n7240), .Y(n5833) );
  NOR2X1 U2722 ( .A(n3482), .B(n5834), .Y(\U3/U94/Z_29 ) );
  NOR2X1 U2723 ( .A(n3482), .B(n5835), .Y(\U3/U94/Z_28 ) );
  NOR2X1 U2724 ( .A(n3482), .B(n5836), .Y(\U3/U94/Z_27 ) );
  NOR2X1 U2725 ( .A(n3482), .B(n5837), .Y(\U3/U94/Z_26 ) );
  NOR2X1 U2726 ( .A(n3482), .B(n5838), .Y(\U3/U94/Z_25 ) );
  NOR2X1 U2727 ( .A(n3482), .B(n5839), .Y(\U3/U94/Z_24 ) );
  NOR2X1 U2728 ( .A(n3482), .B(n5840), .Y(\U3/U94/Z_23 ) );
  NOR2X1 U2729 ( .A(n3482), .B(n5841), .Y(\U3/U94/Z_22 ) );
  NOR2X1 U2730 ( .A(n3482), .B(n5842), .Y(\U3/U94/Z_21 ) );
  NOR2X1 U2731 ( .A(n3482), .B(n5843), .Y(\U3/U94/Z_20 ) );
  OAI21X1 U2732 ( .A(n3844), .B(n5827), .C(n5844), .Y(\U3/U94/Z_2 ) );
  NAND2X1 U2733 ( .A(N2883), .B(n7240), .Y(n5844) );
  NOR2X1 U2734 ( .A(n3482), .B(n5845), .Y(\U3/U94/Z_19 ) );
  NOR2X1 U2735 ( .A(n3482), .B(n5846), .Y(\U3/U94/Z_18 ) );
  NOR2X1 U2736 ( .A(n3482), .B(n5847), .Y(\U3/U94/Z_17 ) );
  NOR2X1 U2737 ( .A(n3482), .B(n5848), .Y(\U3/U94/Z_16 ) );
  NOR2X1 U2738 ( .A(n3482), .B(n5849), .Y(\U3/U94/Z_15 ) );
  NOR2X1 U2739 ( .A(n3482), .B(n5850), .Y(\U3/U94/Z_14 ) );
  AND2X1 U2740 ( .A(N2894), .B(n7240), .Y(\U3/U94/Z_13 ) );
  AND2X1 U2741 ( .A(N2893), .B(n7240), .Y(\U3/U94/Z_12 ) );
  AND2X1 U2742 ( .A(N2892), .B(n7240), .Y(\U3/U94/Z_11 ) );
  AND2X1 U2743 ( .A(N2891), .B(n7240), .Y(\U3/U94/Z_10 ) );
  OAI21X1 U2744 ( .A(n3843), .B(n5827), .C(n5851), .Y(\U3/U94/Z_1 ) );
  NAND2X1 U2745 ( .A(N2882), .B(n7240), .Y(n5851) );
  OAI21X1 U2746 ( .A(n3841), .B(n5827), .C(n5852), .Y(\U3/U94/Z_0 ) );
  NAND2X1 U2747 ( .A(N2881), .B(n7240), .Y(n5852) );
  OAI21X1 U2748 ( .A(n3481), .B(n5744), .C(n3494), .Y(\U3/U93/Z_9 ) );
  NAND2X1 U2749 ( .A(fGy[9]), .B(n7240), .Y(n3494) );
  OAI21X1 U2750 ( .A(n3481), .B(n5742), .C(n3495), .Y(\U3/U93/Z_8 ) );
  NAND2X1 U2751 ( .A(fGy[8]), .B(n7240), .Y(n3495) );
  OAI21X1 U2752 ( .A(n3481), .B(n5740), .C(n5853), .Y(\U3/U93/Z_7 ) );
  AOI21X1 U2753 ( .A(n7246), .B(n5854), .C(\U3/U121/Z_7 ), .Y(n5853) );
  NAND3X1 U2754 ( .A(n5855), .B(n5856), .C(n5857), .Y(n5854) );
  NOR2X1 U2755 ( .A(n5858), .B(n5859), .Y(n5857) );
  OR2X1 U2756 ( .A(n5860), .B(n5861), .Y(n5859) );
  OAI21X1 U2757 ( .A(n3784), .B(n5862), .C(n5863), .Y(n5861) );
  AOI22X1 U2758 ( .A(n5864), .B(\regX[16][7] ), .C(n5865), .D(\regX[20][7] ), 
        .Y(n5863) );
  OAI21X1 U2759 ( .A(n3767), .B(n5866), .C(n5867), .Y(n5860) );
  AOI22X1 U2760 ( .A(n5868), .B(N1742), .C(n5869), .D(\regX[19][7] ), .Y(n5867) );
  INVX1 U2761 ( .A(\regX[13][7] ), .Y(n3767) );
  NAND3X1 U2762 ( .A(n5870), .B(n5871), .C(n5872), .Y(n5858) );
  AOI21X1 U2763 ( .A(n5873), .B(\regX[15][7] ), .C(n5874), .Y(n5872) );
  OAI22X1 U2764 ( .A(n3575), .B(n5875), .C(n3595), .D(n5876), .Y(n5874) );
  AOI22X1 U2765 ( .A(n5877), .B(\regX[18][7] ), .C(n5878), .D(\regX[21][7] ), 
        .Y(n5871) );
  AOI22X1 U2766 ( .A(n5879), .B(\regX[22][7] ), .C(n5880), .D(\regX[17][7] ), 
        .Y(n5870) );
  NOR2X1 U2767 ( .A(n5881), .B(n5882), .Y(n5856) );
  OAI21X1 U2768 ( .A(n3849), .B(n5883), .C(n5884), .Y(n5882) );
  AOI22X1 U2769 ( .A(n5885), .B(\regX[8][7] ), .C(n5886), .D(\regX[7][7] ), 
        .Y(n5884) );
  OAI21X1 U2770 ( .A(n3813), .B(n5887), .C(n5888), .Y(n5881) );
  AOI22X1 U2771 ( .A(n5889), .B(\regX[11][7] ), .C(n5890), .D(N1622), .Y(n5888) );
  NOR2X1 U2772 ( .A(n5891), .B(n5892), .Y(n5855) );
  OAI21X1 U2773 ( .A(n3932), .B(n5893), .C(n5894), .Y(n5892) );
  AOI22X1 U2774 ( .A(n5895), .B(N1382), .C(n5896), .D(\regX[1][7] ), .Y(n5894)
         );
  OAI21X1 U2775 ( .A(n3899), .B(n5897), .C(n5898), .Y(n5891) );
  AOI22X1 U2776 ( .A(n5899), .B(\regX[5][7] ), .C(n5900), .D(N1440), .Y(n5898)
         );
  OAI21X1 U2777 ( .A(n3481), .B(n5738), .C(n5901), .Y(\U3/U93/Z_6 ) );
  AOI21X1 U2778 ( .A(n7246), .B(n5902), .C(\U3/U121/Z_6 ), .Y(n5901) );
  NAND3X1 U2779 ( .A(n5903), .B(n5904), .C(n5905), .Y(n5902) );
  NOR2X1 U2780 ( .A(n5906), .B(n5907), .Y(n5905) );
  OR2X1 U2781 ( .A(n5908), .B(n5909), .Y(n5907) );
  OAI21X1 U2782 ( .A(n3783), .B(n5862), .C(n5910), .Y(n5909) );
  AOI22X1 U2783 ( .A(n5864), .B(\regX[16][6] ), .C(n5865), .D(\regX[20][6] ), 
        .Y(n5910) );
  OAI21X1 U2784 ( .A(n3775), .B(n5866), .C(n5911), .Y(n5908) );
  AOI22X1 U2785 ( .A(n5868), .B(N1741), .C(n5869), .D(\regX[19][6] ), .Y(n5911) );
  INVX1 U2786 ( .A(\regX[13][6] ), .Y(n3775) );
  NAND3X1 U2787 ( .A(n5912), .B(n5913), .C(n5914), .Y(n5906) );
  AOI21X1 U2788 ( .A(n5873), .B(\regX[15][6] ), .C(n5915), .Y(n5914) );
  OAI22X1 U2789 ( .A(n3573), .B(n5875), .C(n3594), .D(n5876), .Y(n5915) );
  AOI22X1 U2790 ( .A(n5877), .B(\regX[18][6] ), .C(n5878), .D(\regX[21][6] ), 
        .Y(n5913) );
  AOI22X1 U2791 ( .A(n5879), .B(\regX[22][6] ), .C(n5880), .D(\regX[17][6] ), 
        .Y(n5912) );
  NOR2X1 U2792 ( .A(n5916), .B(n5917), .Y(n5904) );
  OAI21X1 U2793 ( .A(n3848), .B(n5883), .C(n5918), .Y(n5917) );
  AOI22X1 U2794 ( .A(n5885), .B(\regX[8][6] ), .C(n5886), .D(\regX[7][6] ), 
        .Y(n5918) );
  OAI21X1 U2795 ( .A(n3812), .B(n5887), .C(n5919), .Y(n5916) );
  AOI22X1 U2796 ( .A(n5889), .B(\regX[11][6] ), .C(n5890), .D(N1621), .Y(n5919) );
  NOR2X1 U2797 ( .A(n5920), .B(n5921), .Y(n5903) );
  OAI21X1 U2798 ( .A(n3931), .B(n5893), .C(n5922), .Y(n5921) );
  AOI22X1 U2799 ( .A(n5895), .B(N1381), .C(n5896), .D(\regX[1][6] ), .Y(n5922)
         );
  OAI21X1 U2800 ( .A(n3898), .B(n5897), .C(n5923), .Y(n5920) );
  AOI22X1 U2801 ( .A(n5899), .B(\regX[5][6] ), .C(n5900), .D(N1439), .Y(n5923)
         );
  OAI21X1 U2802 ( .A(n3481), .B(n5736), .C(n5924), .Y(\U3/U93/Z_5 ) );
  AOI21X1 U2803 ( .A(n7246), .B(n5925), .C(\U3/U121/Z_5 ), .Y(n5924) );
  NAND3X1 U2804 ( .A(n5926), .B(n5927), .C(n5928), .Y(n5925) );
  NOR2X1 U2805 ( .A(n5929), .B(n5930), .Y(n5928) );
  OR2X1 U2806 ( .A(n5931), .B(n5932), .Y(n5930) );
  OAI21X1 U2807 ( .A(n3782), .B(n5862), .C(n5933), .Y(n5932) );
  AOI22X1 U2808 ( .A(n5864), .B(\regX[16][5] ), .C(n5865), .D(\regX[20][5] ), 
        .Y(n5933) );
  OAI21X1 U2809 ( .A(n3774), .B(n5866), .C(n5934), .Y(n5931) );
  AOI22X1 U2810 ( .A(n5868), .B(N1740), .C(n5869), .D(\regX[19][5] ), .Y(n5934) );
  INVX1 U2811 ( .A(\regX[13][5] ), .Y(n3774) );
  NAND3X1 U2812 ( .A(n5935), .B(n5936), .C(n5937), .Y(n5929) );
  AOI21X1 U2813 ( .A(n5873), .B(\regX[15][5] ), .C(n5938), .Y(n5937) );
  OAI22X1 U2814 ( .A(n3571), .B(n5875), .C(n3593), .D(n5876), .Y(n5938) );
  AOI22X1 U2815 ( .A(n5877), .B(\regX[18][5] ), .C(n5878), .D(\regX[21][5] ), 
        .Y(n5936) );
  AOI22X1 U2816 ( .A(n5879), .B(\regX[22][5] ), .C(n5880), .D(\regX[17][5] ), 
        .Y(n5935) );
  NOR2X1 U2817 ( .A(n5939), .B(n5940), .Y(n5927) );
  OAI21X1 U2818 ( .A(n3847), .B(n5883), .C(n5941), .Y(n5940) );
  AOI22X1 U2819 ( .A(n5885), .B(\regX[8][5] ), .C(n5886), .D(\regX[7][5] ), 
        .Y(n5941) );
  OAI21X1 U2820 ( .A(n3811), .B(n5887), .C(n5942), .Y(n5939) );
  AOI22X1 U2821 ( .A(n5889), .B(\regX[11][5] ), .C(n5890), .D(N1620), .Y(n5942) );
  NOR2X1 U2822 ( .A(n5943), .B(n5944), .Y(n5926) );
  OAI21X1 U2823 ( .A(n3930), .B(n5893), .C(n5945), .Y(n5944) );
  AOI22X1 U2824 ( .A(n5895), .B(N1380), .C(n5896), .D(\regX[1][5] ), .Y(n5945)
         );
  OAI21X1 U2825 ( .A(n3897), .B(n5897), .C(n5946), .Y(n5943) );
  AOI22X1 U2826 ( .A(n5899), .B(\regX[5][5] ), .C(n5900), .D(N1438), .Y(n5946)
         );
  OAI21X1 U2827 ( .A(n3481), .B(n5734), .C(n5947), .Y(\U3/U93/Z_4 ) );
  AOI21X1 U2828 ( .A(n7246), .B(n5948), .C(\U3/U121/Z_4 ), .Y(n5947) );
  NAND3X1 U2829 ( .A(n5949), .B(n5950), .C(n5951), .Y(n5948) );
  NOR2X1 U2830 ( .A(n5952), .B(n5953), .Y(n5951) );
  OR2X1 U2831 ( .A(n5954), .B(n5955), .Y(n5953) );
  OAI21X1 U2832 ( .A(n3781), .B(n5862), .C(n5956), .Y(n5955) );
  AOI22X1 U2833 ( .A(n5864), .B(\regX[16][4] ), .C(n5865), .D(\regX[20][4] ), 
        .Y(n5956) );
  OAI21X1 U2834 ( .A(n3773), .B(n5866), .C(n5957), .Y(n5954) );
  AOI22X1 U2835 ( .A(n5868), .B(N1739), .C(n5869), .D(\regX[19][4] ), .Y(n5957) );
  INVX1 U2836 ( .A(\regX[13][4] ), .Y(n3773) );
  NAND3X1 U2837 ( .A(n5958), .B(n5959), .C(n5960), .Y(n5952) );
  AOI21X1 U2838 ( .A(n5873), .B(\regX[15][4] ), .C(n5961), .Y(n5960) );
  OAI22X1 U2839 ( .A(n3569), .B(n5875), .C(n3592), .D(n5876), .Y(n5961) );
  AOI22X1 U2840 ( .A(n5877), .B(\regX[18][4] ), .C(n5878), .D(\regX[21][4] ), 
        .Y(n5959) );
  AOI22X1 U2841 ( .A(n5879), .B(\regX[22][4] ), .C(n5880), .D(\regX[17][4] ), 
        .Y(n5958) );
  NOR2X1 U2842 ( .A(n5962), .B(n5963), .Y(n5950) );
  OAI21X1 U2843 ( .A(n3846), .B(n5883), .C(n5964), .Y(n5963) );
  AOI22X1 U2844 ( .A(n5885), .B(\regX[8][4] ), .C(n5886), .D(\regX[7][4] ), 
        .Y(n5964) );
  OAI21X1 U2845 ( .A(n3810), .B(n5887), .C(n5965), .Y(n5962) );
  AOI22X1 U2846 ( .A(n5889), .B(\regX[11][4] ), .C(n5890), .D(N1619), .Y(n5965) );
  NOR2X1 U2847 ( .A(n5966), .B(n5967), .Y(n5949) );
  OAI21X1 U2848 ( .A(n3929), .B(n5893), .C(n5968), .Y(n5967) );
  AOI22X1 U2849 ( .A(n5895), .B(N1379), .C(n5896), .D(\regX[1][4] ), .Y(n5968)
         );
  OAI21X1 U2850 ( .A(n3896), .B(n5897), .C(n5969), .Y(n5966) );
  AOI22X1 U2851 ( .A(n5899), .B(\regX[5][4] ), .C(n5900), .D(N1437), .Y(n5969)
         );
  OAI21X1 U2852 ( .A(n3481), .B(n5788), .C(n3496), .Y(\U3/U93/Z_31 ) );
  NAND2X1 U2853 ( .A(n7240), .B(fGy[31]), .Y(n3496) );
  OAI21X1 U2854 ( .A(n3481), .B(n5786), .C(n3497), .Y(\U3/U93/Z_30 ) );
  NAND2X1 U2855 ( .A(fGy[30]), .B(n7240), .Y(n3497) );
  OAI21X1 U2856 ( .A(n3481), .B(n5732), .C(n5970), .Y(\U3/U93/Z_3 ) );
  AOI22X1 U2857 ( .A(n7246), .B(n5971), .C(fGy[3]), .D(n7240), .Y(n5970) );
  NAND3X1 U2858 ( .A(n5972), .B(n5973), .C(n5974), .Y(n5971) );
  NOR2X1 U2859 ( .A(n5975), .B(n5976), .Y(n5974) );
  OR2X1 U2860 ( .A(n5977), .B(n5978), .Y(n5976) );
  OAI21X1 U2861 ( .A(n3780), .B(n5862), .C(n5979), .Y(n5978) );
  AOI22X1 U2862 ( .A(n5864), .B(\regX[16][3] ), .C(n5865), .D(\regX[20][3] ), 
        .Y(n5979) );
  OAI21X1 U2863 ( .A(n3772), .B(n5866), .C(n5980), .Y(n5977) );
  AOI22X1 U2864 ( .A(n5868), .B(N1738), .C(n5869), .D(\regX[19][3] ), .Y(n5980) );
  INVX1 U2865 ( .A(\regX[13][3] ), .Y(n3772) );
  NAND3X1 U2866 ( .A(n5981), .B(n5982), .C(n5983), .Y(n5975) );
  AOI21X1 U2867 ( .A(n5873), .B(\regX[15][3] ), .C(n5984), .Y(n5983) );
  OAI22X1 U2868 ( .A(n3567), .B(n5875), .C(n3591), .D(n5876), .Y(n5984) );
  AOI22X1 U2869 ( .A(n5877), .B(\regX[18][3] ), .C(n5878), .D(\regX[21][3] ), 
        .Y(n5982) );
  AOI22X1 U2870 ( .A(n5879), .B(\regX[22][3] ), .C(n5880), .D(\regX[17][3] ), 
        .Y(n5981) );
  NOR2X1 U2871 ( .A(n5985), .B(n5986), .Y(n5973) );
  OAI21X1 U2872 ( .A(n3845), .B(n5883), .C(n5987), .Y(n5986) );
  AOI22X1 U2873 ( .A(n5885), .B(\regX[8][3] ), .C(n5886), .D(\regX[7][3] ), 
        .Y(n5987) );
  OAI21X1 U2874 ( .A(n3809), .B(n5887), .C(n5988), .Y(n5985) );
  AOI22X1 U2875 ( .A(n5889), .B(\regX[11][3] ), .C(n5890), .D(N1618), .Y(n5988) );
  NOR2X1 U2876 ( .A(n5989), .B(n5990), .Y(n5972) );
  OAI21X1 U2877 ( .A(n3928), .B(n5893), .C(n5991), .Y(n5990) );
  AOI22X1 U2878 ( .A(n5895), .B(N1378), .C(n5896), .D(\regX[1][3] ), .Y(n5991)
         );
  OAI21X1 U2879 ( .A(n3895), .B(n5897), .C(n5992), .Y(n5989) );
  AOI22X1 U2880 ( .A(n5899), .B(\regX[5][3] ), .C(n5900), .D(N1436), .Y(n5992)
         );
  OAI21X1 U2881 ( .A(n3481), .B(n5784), .C(n3498), .Y(\U3/U93/Z_29 ) );
  NAND2X1 U2882 ( .A(fGy[29]), .B(n7240), .Y(n3498) );
  OAI21X1 U2883 ( .A(n3481), .B(n5782), .C(n3499), .Y(\U3/U93/Z_28 ) );
  NAND2X1 U2884 ( .A(fGy[28]), .B(n7240), .Y(n3499) );
  OAI21X1 U2885 ( .A(n3481), .B(n5780), .C(n3500), .Y(\U3/U93/Z_27 ) );
  NAND2X1 U2886 ( .A(fGy[27]), .B(n7240), .Y(n3500) );
  OAI21X1 U2887 ( .A(n3481), .B(n5778), .C(n3501), .Y(\U3/U93/Z_26 ) );
  NAND2X1 U2888 ( .A(fGy[26]), .B(n7240), .Y(n3501) );
  OAI21X1 U2889 ( .A(n3481), .B(n5776), .C(n3502), .Y(\U3/U93/Z_25 ) );
  NAND2X1 U2890 ( .A(fGy[25]), .B(n7240), .Y(n3502) );
  OAI21X1 U2891 ( .A(n3481), .B(n5774), .C(n3503), .Y(\U3/U93/Z_24 ) );
  NAND2X1 U2892 ( .A(fGy[24]), .B(n7240), .Y(n3503) );
  OAI21X1 U2893 ( .A(n3481), .B(n5772), .C(n3504), .Y(\U3/U93/Z_23 ) );
  NAND2X1 U2894 ( .A(fGy[23]), .B(n7240), .Y(n3504) );
  OAI21X1 U2895 ( .A(n3481), .B(n5770), .C(n3505), .Y(\U3/U93/Z_22 ) );
  NAND2X1 U2896 ( .A(fGy[22]), .B(n7240), .Y(n3505) );
  OAI21X1 U2897 ( .A(n3481), .B(n5768), .C(n3506), .Y(\U3/U93/Z_21 ) );
  NAND2X1 U2898 ( .A(fGy[21]), .B(n7240), .Y(n3506) );
  OAI21X1 U2899 ( .A(n3481), .B(n5766), .C(n3507), .Y(\U3/U93/Z_20 ) );
  NAND2X1 U2900 ( .A(fGy[20]), .B(n7240), .Y(n3507) );
  OAI21X1 U2901 ( .A(n3481), .B(n5730), .C(n5993), .Y(\U3/U93/Z_2 ) );
  AOI22X1 U2902 ( .A(n7246), .B(n5994), .C(fGy[2]), .D(n7240), .Y(n5993) );
  NAND3X1 U2903 ( .A(n5995), .B(n5996), .C(n5997), .Y(n5994) );
  NOR2X1 U2904 ( .A(n5998), .B(n5999), .Y(n5997) );
  OR2X1 U2905 ( .A(n6000), .B(n6001), .Y(n5999) );
  OAI21X1 U2906 ( .A(n3779), .B(n5862), .C(n6002), .Y(n6001) );
  AOI22X1 U2907 ( .A(n5864), .B(\regX[16][2] ), .C(n5865), .D(\regX[20][2] ), 
        .Y(n6002) );
  OAI21X1 U2908 ( .A(n3771), .B(n5866), .C(n6003), .Y(n6000) );
  AOI22X1 U2909 ( .A(n5868), .B(N1737), .C(n5869), .D(\regX[19][2] ), .Y(n6003) );
  INVX1 U2910 ( .A(\regX[13][2] ), .Y(n3771) );
  NAND3X1 U2911 ( .A(n6004), .B(n6005), .C(n6006), .Y(n5998) );
  AOI21X1 U2912 ( .A(n5873), .B(\regX[15][2] ), .C(n6007), .Y(n6006) );
  OAI22X1 U2913 ( .A(n3565), .B(n5875), .C(n3590), .D(n5876), .Y(n6007) );
  AOI22X1 U2914 ( .A(n5877), .B(\regX[18][2] ), .C(n5878), .D(\regX[21][2] ), 
        .Y(n6005) );
  AOI22X1 U2915 ( .A(n5879), .B(\regX[22][2] ), .C(n5880), .D(\regX[17][2] ), 
        .Y(n6004) );
  NOR2X1 U2916 ( .A(n6008), .B(n6009), .Y(n5996) );
  OAI21X1 U2917 ( .A(n3844), .B(n5883), .C(n6010), .Y(n6009) );
  AOI22X1 U2918 ( .A(n5885), .B(\regX[8][2] ), .C(n5886), .D(\regX[7][2] ), 
        .Y(n6010) );
  OAI21X1 U2919 ( .A(n3808), .B(n5887), .C(n6011), .Y(n6008) );
  AOI22X1 U2920 ( .A(n5889), .B(\regX[11][2] ), .C(n5890), .D(N1617), .Y(n6011) );
  NOR2X1 U2921 ( .A(n6012), .B(n6013), .Y(n5995) );
  OAI21X1 U2922 ( .A(n3926), .B(n5893), .C(n6014), .Y(n6013) );
  AOI22X1 U2923 ( .A(n5895), .B(N1377), .C(n5896), .D(\regX[1][2] ), .Y(n6014)
         );
  OAI21X1 U2924 ( .A(n3894), .B(n5897), .C(n6015), .Y(n6012) );
  AOI22X1 U2925 ( .A(n5899), .B(\regX[5][2] ), .C(n5900), .D(N1435), .Y(n6015)
         );
  OAI21X1 U2926 ( .A(n3481), .B(n5764), .C(n3508), .Y(\U3/U93/Z_19 ) );
  NAND2X1 U2927 ( .A(fGy[19]), .B(n7240), .Y(n3508) );
  OAI21X1 U2928 ( .A(n3481), .B(n5762), .C(n3509), .Y(\U3/U93/Z_18 ) );
  NAND2X1 U2929 ( .A(fGy[18]), .B(n7240), .Y(n3509) );
  OAI21X1 U2930 ( .A(n3481), .B(n5760), .C(n3510), .Y(\U3/U93/Z_17 ) );
  NAND2X1 U2931 ( .A(fGy[17]), .B(n7240), .Y(n3510) );
  OAI21X1 U2932 ( .A(n3481), .B(n5758), .C(n3511), .Y(\U3/U93/Z_16 ) );
  NAND2X1 U2933 ( .A(fGy[16]), .B(n7240), .Y(n3511) );
  OAI21X1 U2934 ( .A(n3481), .B(n5756), .C(n3512), .Y(\U3/U93/Z_15 ) );
  NAND2X1 U2935 ( .A(fGy[15]), .B(n7240), .Y(n3512) );
  OAI21X1 U2936 ( .A(n3481), .B(n5754), .C(n3513), .Y(\U3/U93/Z_14 ) );
  NAND2X1 U2937 ( .A(fGy[14]), .B(n7240), .Y(n3513) );
  OAI21X1 U2938 ( .A(n3481), .B(n5752), .C(n3514), .Y(\U3/U93/Z_13 ) );
  NAND2X1 U2939 ( .A(fGy[13]), .B(n7240), .Y(n3514) );
  OAI21X1 U2940 ( .A(n3481), .B(n5750), .C(n3515), .Y(\U3/U93/Z_12 ) );
  NAND2X1 U2941 ( .A(fGy[12]), .B(n7240), .Y(n3515) );
  OAI21X1 U2942 ( .A(n3481), .B(n5748), .C(n3516), .Y(\U3/U93/Z_11 ) );
  NAND2X1 U2943 ( .A(fGy[11]), .B(n7240), .Y(n3516) );
  OAI21X1 U2944 ( .A(n3481), .B(n5746), .C(n3517), .Y(\U3/U93/Z_10 ) );
  NAND2X1 U2945 ( .A(fGy[10]), .B(n7240), .Y(n3517) );
  OAI21X1 U2946 ( .A(n3481), .B(n5728), .C(n6016), .Y(\U3/U93/Z_1 ) );
  AOI22X1 U2947 ( .A(n7246), .B(n6017), .C(fGy[1]), .D(n7240), .Y(n6016) );
  NAND3X1 U2948 ( .A(n6018), .B(n6019), .C(n6020), .Y(n6017) );
  NOR2X1 U2949 ( .A(n6021), .B(n6022), .Y(n6020) );
  OR2X1 U2950 ( .A(n6023), .B(n6024), .Y(n6022) );
  OAI21X1 U2951 ( .A(n3778), .B(n5862), .C(n6025), .Y(n6024) );
  AOI22X1 U2952 ( .A(n5864), .B(\regX[16][1] ), .C(n5865), .D(\regX[20][1] ), 
        .Y(n6025) );
  OAI21X1 U2953 ( .A(n3770), .B(n5866), .C(n6026), .Y(n6023) );
  AOI22X1 U2954 ( .A(n5868), .B(N1736), .C(n5869), .D(\regX[19][1] ), .Y(n6026) );
  INVX1 U2955 ( .A(\regX[13][1] ), .Y(n3770) );
  NAND3X1 U2956 ( .A(n6027), .B(n6028), .C(n6029), .Y(n6021) );
  AOI21X1 U2957 ( .A(n5873), .B(\regX[15][1] ), .C(n6030), .Y(n6029) );
  OAI22X1 U2958 ( .A(n3563), .B(n5875), .C(n3589), .D(n5876), .Y(n6030) );
  AOI22X1 U2959 ( .A(n5877), .B(\regX[18][1] ), .C(n5878), .D(\regX[21][1] ), 
        .Y(n6028) );
  AOI22X1 U2960 ( .A(n5879), .B(\regX[22][1] ), .C(n5880), .D(\regX[17][1] ), 
        .Y(n6027) );
  NOR2X1 U2961 ( .A(n6031), .B(n6032), .Y(n6019) );
  OAI21X1 U2962 ( .A(n3843), .B(n5883), .C(n6033), .Y(n6032) );
  AOI22X1 U2963 ( .A(n5885), .B(\regX[8][1] ), .C(n5886), .D(\regX[7][1] ), 
        .Y(n6033) );
  OAI21X1 U2964 ( .A(n3807), .B(n5887), .C(n6034), .Y(n6031) );
  AOI22X1 U2965 ( .A(n5889), .B(\regX[11][1] ), .C(n5890), .D(N1616), .Y(n6034) );
  NOR2X1 U2966 ( .A(n6035), .B(n6036), .Y(n6018) );
  OAI21X1 U2967 ( .A(n3934), .B(n5893), .C(n6037), .Y(n6036) );
  AOI22X1 U2968 ( .A(n5895), .B(N1376), .C(n5896), .D(\regX[1][1] ), .Y(n6037)
         );
  OAI21X1 U2969 ( .A(n3893), .B(n5897), .C(n6038), .Y(n6035) );
  AOI22X1 U2970 ( .A(n5899), .B(\regX[5][1] ), .C(n5900), .D(N1434), .Y(n6038)
         );
  OAI21X1 U2971 ( .A(n3481), .B(n5726), .C(n6039), .Y(\U3/U93/Z_0 ) );
  AOI22X1 U2972 ( .A(n7246), .B(n6040), .C(fGy[0]), .D(n7240), .Y(n6039) );
  NAND3X1 U2973 ( .A(n6041), .B(n6042), .C(n6043), .Y(n6040) );
  NOR2X1 U2974 ( .A(n6044), .B(n6045), .Y(n6043) );
  OR2X1 U2975 ( .A(n6046), .B(n6047), .Y(n6045) );
  OAI21X1 U2976 ( .A(n3776), .B(n5862), .C(n6048), .Y(n6047) );
  AOI22X1 U2977 ( .A(n5864), .B(\regX[16][0] ), .C(n5865), .D(\regX[20][0] ), 
        .Y(n6048) );
  AND2X1 U2978 ( .A(n6049), .B(n6050), .Y(n5865) );
  INVX1 U2979 ( .A(n6051), .Y(n5864) );
  NAND3X1 U2980 ( .A(n6050), .B(n6052), .C(n6053), .Y(n6051) );
  NAND2X1 U2981 ( .A(n6054), .B(n6049), .Y(n5862) );
  OAI21X1 U2982 ( .A(n3769), .B(n5866), .C(n6055), .Y(n6046) );
  AOI22X1 U2983 ( .A(n5868), .B(N1735), .C(n5869), .D(\regX[19][0] ), .Y(n6055) );
  AND2X1 U2984 ( .A(n6056), .B(n6057), .Y(n5869) );
  AND2X1 U2985 ( .A(n6054), .B(n6058), .Y(n5868) );
  NAND2X1 U2986 ( .A(n6059), .B(n6049), .Y(n5866) );
  INVX1 U2987 ( .A(\regX[13][0] ), .Y(n3769) );
  NAND3X1 U2988 ( .A(n6060), .B(n6061), .C(n6062), .Y(n6044) );
  AOI21X1 U2989 ( .A(n5873), .B(\regX[15][0] ), .C(n6063), .Y(n6062) );
  OAI22X1 U2990 ( .A(n3560), .B(n5875), .C(n3587), .D(n5876), .Y(n6063) );
  NAND2X1 U2991 ( .A(n6058), .B(n6056), .Y(n5876) );
  NAND2X1 U2992 ( .A(n6064), .B(n6065), .Y(n5875) );
  INVX1 U2993 ( .A(n6066), .Y(n6065) );
  AND2X1 U2994 ( .A(n6059), .B(n6058), .Y(n5873) );
  AOI22X1 U2995 ( .A(n5877), .B(\regX[18][0] ), .C(n5878), .D(\regX[21][0] ), 
        .Y(n6061) );
  AND2X1 U2996 ( .A(n6049), .B(n6056), .Y(n5878) );
  AND2X1 U2997 ( .A(n6057), .B(n6050), .Y(n5877) );
  AOI22X1 U2998 ( .A(n5879), .B(\regX[22][0] ), .C(n5880), .D(\regX[17][0] ), 
        .Y(n6060) );
  AND2X1 U2999 ( .A(n6053), .B(n6056), .Y(n5880) );
  NOR2X1 U3000 ( .A(n6066), .B(n6067), .Y(n6056) );
  AND2X1 U3001 ( .A(n6058), .B(n6050), .Y(n5879) );
  NOR2X1 U3002 ( .A(n6068), .B(n6066), .Y(n6050) );
  NOR2X1 U3003 ( .A(n6069), .B(n6070), .Y(n6042) );
  OAI21X1 U3004 ( .A(n3841), .B(n5883), .C(n6071), .Y(n6070) );
  AOI22X1 U3005 ( .A(n5885), .B(\regX[8][0] ), .C(n5886), .D(\regX[7][0] ), 
        .Y(n6071) );
  AND2X1 U3006 ( .A(n6072), .B(n6058), .Y(n5886) );
  INVX1 U3007 ( .A(n6073), .Y(n5885) );
  NAND3X1 U3008 ( .A(n6053), .B(n6066), .C(n6054), .Y(n6073) );
  NAND2X1 U3009 ( .A(n6074), .B(n6058), .Y(n5883) );
  NOR2X1 U3010 ( .A(n6075), .B(n6076), .Y(n6058) );
  OAI21X1 U3011 ( .A(n3805), .B(n5887), .C(n6077), .Y(n6069) );
  AOI22X1 U3012 ( .A(n5889), .B(\regX[11][0] ), .C(n5890), .D(N1615), .Y(n6077) );
  AND2X1 U3013 ( .A(n6054), .B(n6057), .Y(n5890) );
  NOR2X1 U3014 ( .A(n6052), .B(n6068), .Y(n6054) );
  AND2X1 U3015 ( .A(n6059), .B(n6057), .Y(n5889) );
  NAND2X1 U3016 ( .A(n6059), .B(n6053), .Y(n5887) );
  NOR2X1 U3017 ( .A(n6052), .B(n6067), .Y(n6059) );
  NOR2X1 U3018 ( .A(n6078), .B(n6079), .Y(n6041) );
  OAI21X1 U3019 ( .A(n3933), .B(n5893), .C(n6080), .Y(n6079) );
  AOI22X1 U3020 ( .A(n5895), .B(N1375), .C(n5896), .D(\regX[1][0] ), .Y(n6080)
         );
  AND2X1 U3021 ( .A(n6072), .B(n6053), .Y(n5896) );
  AND2X1 U3022 ( .A(n6074), .B(n6057), .Y(n5895) );
  NAND2X1 U3023 ( .A(n6074), .B(n6053), .Y(n5893) );
  NOR2X1 U3024 ( .A(n6081), .B(n6082), .Y(n6053) );
  OAI21X1 U3025 ( .A(n3891), .B(n5897), .C(n6083), .Y(n6078) );
  AOI22X1 U3026 ( .A(n5899), .B(\regX[5][0] ), .C(n5900), .D(N1433), .Y(n6083)
         );
  AND2X1 U3027 ( .A(n6074), .B(n6049), .Y(n5900) );
  INVX1 U3028 ( .A(n6084), .Y(n6074) );
  NAND3X1 U3029 ( .A(n6052), .B(n6066), .C(n6067), .Y(n6084) );
  INVX1 U3030 ( .A(n6068), .Y(n6067) );
  AND2X1 U3031 ( .A(n6072), .B(n6049), .Y(n5899) );
  NOR2X1 U3032 ( .A(n6081), .B(n6075), .Y(n6049) );
  NAND2X1 U3033 ( .A(n6072), .B(n6057), .Y(n5897) );
  NOR2X1 U3034 ( .A(n6082), .B(n6076), .Y(n6057) );
  INVX1 U3035 ( .A(n6085), .Y(n6072) );
  NAND3X1 U3036 ( .A(n6066), .B(n6068), .C(n6052), .Y(n6085) );
  INVX1 U3037 ( .A(n6064), .Y(n6052) );
  OAI21X1 U3038 ( .A(n3475), .B(n3630), .C(n6086), .Y(\U3/U91/Z_7 ) );
  OAI21X1 U3039 ( .A(n3475), .B(n3629), .C(n6086), .Y(\U3/U91/Z_6 ) );
  OAI21X1 U3040 ( .A(n3475), .B(n3628), .C(n6086), .Y(\U3/U91/Z_5 ) );
  OAI21X1 U3041 ( .A(n3475), .B(n3627), .C(n6086), .Y(\U3/U91/Z_4 ) );
  OAI21X1 U3042 ( .A(n3475), .B(n3626), .C(n6086), .Y(\U3/U91/Z_3 ) );
  OAI21X1 U3043 ( .A(n3475), .B(n3625), .C(n6086), .Y(\U3/U91/Z_2 ) );
  OAI21X1 U3044 ( .A(n3475), .B(n3624), .C(n6086), .Y(\U3/U91/Z_1 ) );
  NAND2X1 U3045 ( .A(dy[1]), .B(n7246), .Y(n6086) );
  OAI22X1 U3046 ( .A(n5827), .B(n5825), .C(n3475), .D(n3622), .Y(\U3/U91/Z_0 )
         );
  NAND2X1 U3047 ( .A(n5827), .B(n3475), .Y(\U3/U90/Z_0 ) );
  OR2X1 U3048 ( .A(\U3/U122/Z_8 ), .B(n3483), .Y(\U3/U88/Z_9 ) );
  OAI21X1 U3049 ( .A(n5826), .B(n4023), .C(n3476), .Y(\U3/U88/Z_8 ) );
  OAI21X1 U3050 ( .A(n3475), .B(n3595), .C(n6087), .Y(\U3/U88/Z_7 ) );
  AOI21X1 U3051 ( .A(fGx[7]), .B(n7240), .C(n3483), .Y(n6087) );
  OAI21X1 U3052 ( .A(n3475), .B(n3594), .C(n6088), .Y(\U3/U88/Z_6 ) );
  AOI21X1 U3053 ( .A(fGx[6]), .B(n7240), .C(n3483), .Y(n6088) );
  OAI21X1 U3054 ( .A(n3475), .B(n3593), .C(n6089), .Y(\U3/U88/Z_5 ) );
  AOI21X1 U3055 ( .A(fGx[5]), .B(n7240), .C(n3483), .Y(n6089) );
  OAI21X1 U3056 ( .A(n3475), .B(n3592), .C(n6090), .Y(\U3/U88/Z_4 ) );
  AOI21X1 U3057 ( .A(fGx[4]), .B(n7240), .C(n3483), .Y(n6090) );
  OR2X1 U3058 ( .A(\U3/U122/Z_29 ), .B(n3483), .Y(\U3/U88/Z_30 ) );
  OAI21X1 U3059 ( .A(n3475), .B(n3591), .C(n6091), .Y(\U3/U88/Z_3 ) );
  AOI21X1 U3060 ( .A(fGx[3]), .B(n7240), .C(n3483), .Y(n6091) );
  OR2X1 U3061 ( .A(\U3/U122/Z_28 ), .B(n3483), .Y(\U3/U88/Z_29 ) );
  OR2X1 U3062 ( .A(\U3/U122/Z_27 ), .B(n3483), .Y(\U3/U88/Z_28 ) );
  OR2X1 U3063 ( .A(\U3/U122/Z_26 ), .B(n3483), .Y(\U3/U88/Z_27 ) );
  OR2X1 U3064 ( .A(\U3/U122/Z_25 ), .B(n3483), .Y(\U3/U88/Z_26 ) );
  OR2X1 U3065 ( .A(\U3/U122/Z_24 ), .B(n3483), .Y(\U3/U88/Z_25 ) );
  OR2X1 U3066 ( .A(\U3/U122/Z_23 ), .B(n3483), .Y(\U3/U88/Z_24 ) );
  OR2X1 U3067 ( .A(\U3/U122/Z_22 ), .B(n3483), .Y(\U3/U88/Z_23 ) );
  OR2X1 U3068 ( .A(\U3/U122/Z_21 ), .B(n3483), .Y(\U3/U88/Z_22 ) );
  OR2X1 U3069 ( .A(\U3/U122/Z_20 ), .B(n3483), .Y(\U3/U88/Z_21 ) );
  OR2X1 U3070 ( .A(\U3/U122/Z_19 ), .B(n3483), .Y(\U3/U88/Z_20 ) );
  OAI21X1 U3071 ( .A(n3475), .B(n3590), .C(n6092), .Y(\U3/U88/Z_2 ) );
  AOI21X1 U3072 ( .A(fGx[2]), .B(n7240), .C(n3483), .Y(n6092) );
  OR2X1 U3073 ( .A(\U3/U122/Z_18 ), .B(n3483), .Y(\U3/U88/Z_19 ) );
  OR2X1 U3074 ( .A(\U3/U122/Z_17 ), .B(n3483), .Y(\U3/U88/Z_18 ) );
  OR2X1 U3075 ( .A(\U3/U122/Z_16 ), .B(n3483), .Y(\U3/U88/Z_17 ) );
  OR2X1 U3076 ( .A(\U3/U122/Z_15 ), .B(n3483), .Y(\U3/U88/Z_16 ) );
  OR2X1 U3077 ( .A(\U3/U122/Z_14 ), .B(n3483), .Y(\U3/U88/Z_15 ) );
  OR2X1 U3078 ( .A(\U3/U122/Z_13 ), .B(n3483), .Y(\U3/U88/Z_14 ) );
  OR2X1 U3079 ( .A(\U3/U122/Z_12 ), .B(n3483), .Y(\U3/U88/Z_13 ) );
  OR2X1 U3080 ( .A(\U3/U122/Z_11 ), .B(n3483), .Y(\U3/U88/Z_12 ) );
  OR2X1 U3081 ( .A(\U3/U122/Z_10 ), .B(n3483), .Y(\U3/U88/Z_11 ) );
  OR2X1 U3082 ( .A(\U3/U122/Z_9 ), .B(n3483), .Y(\U3/U88/Z_10 ) );
  OAI21X1 U3083 ( .A(n3475), .B(n3589), .C(n6093), .Y(\U3/U88/Z_1 ) );
  AOI21X1 U3084 ( .A(fGx[1]), .B(n7240), .C(n3483), .Y(n6093) );
  OAI21X1 U3085 ( .A(n3475), .B(n3587), .C(n6094), .Y(\U3/U88/Z_0 ) );
  AOI21X1 U3086 ( .A(fGx[0]), .B(n7240), .C(n3483), .Y(n6094) );
  NOR2X1 U3087 ( .A(n3476), .B(n3784), .Y(\U3/U87/Z_7 ) );
  NOR2X1 U3088 ( .A(n3476), .B(n3783), .Y(\U3/U87/Z_6 ) );
  NOR2X1 U3089 ( .A(n3476), .B(n3782), .Y(\U3/U87/Z_5 ) );
  NOR2X1 U3090 ( .A(n3476), .B(n3781), .Y(\U3/U87/Z_4 ) );
  NOR2X1 U3091 ( .A(n3476), .B(n3780), .Y(\U3/U87/Z_3 ) );
  OAI21X1 U3092 ( .A(n3476), .B(n3779), .C(n3482), .Y(\U3/U87/Z_2 ) );
  OAI21X1 U3093 ( .A(n3476), .B(n3778), .C(n3475), .Y(\U3/U87/Z_1 ) );
  OAI21X1 U3094 ( .A(n3476), .B(n3776), .C(n6095), .Y(\U3/U87/Z_0 ) );
  NOR2X1 U3095 ( .A(n7253), .B(n7240), .Y(n6095) );
  OAI21X1 U3096 ( .A(n3477), .B(n4026), .C(n3476), .Y(\U3/U85/Z_9 ) );
  OAI21X1 U3097 ( .A(n3477), .B(n4023), .C(n3476), .Y(\U3/U85/Z_8 ) );
  OAI21X1 U3098 ( .A(n3477), .B(n6096), .C(n6097), .Y(\U3/U85/Z_7 ) );
  AOI21X1 U3099 ( .A(\regX[22][7] ), .B(n7253), .C(n3483), .Y(n6097) );
  OAI21X1 U3100 ( .A(n3477), .B(n6098), .C(n6099), .Y(\U3/U85/Z_6 ) );
  AOI21X1 U3101 ( .A(\regX[22][6] ), .B(n7253), .C(n3483), .Y(n6099) );
  OAI21X1 U3102 ( .A(n3477), .B(n6100), .C(n6101), .Y(\U3/U85/Z_5 ) );
  AOI21X1 U3103 ( .A(\regX[22][5] ), .B(n7253), .C(n3483), .Y(n6101) );
  OAI21X1 U3104 ( .A(n3477), .B(n6102), .C(n6103), .Y(\U3/U85/Z_4 ) );
  AOI21X1 U3105 ( .A(\regX[22][4] ), .B(n7253), .C(n3483), .Y(n6103) );
  OAI21X1 U3106 ( .A(n3477), .B(n4070), .C(n3476), .Y(\U3/U85/Z_31 ) );
  OAI21X1 U3107 ( .A(n3477), .B(n4068), .C(n3476), .Y(\U3/U85/Z_30 ) );
  OAI21X1 U3108 ( .A(n3477), .B(n6104), .C(n6105), .Y(\U3/U85/Z_3 ) );
  AOI21X1 U3109 ( .A(\regX[22][3] ), .B(n7253), .C(n3483), .Y(n6105) );
  OAI21X1 U3110 ( .A(n3477), .B(n4066), .C(n3476), .Y(\U3/U85/Z_29 ) );
  OAI21X1 U3111 ( .A(n3477), .B(n4064), .C(n3476), .Y(\U3/U85/Z_28 ) );
  OAI21X1 U3112 ( .A(n3477), .B(n4062), .C(n3476), .Y(\U3/U85/Z_27 ) );
  OAI21X1 U3113 ( .A(n3477), .B(n4060), .C(n3476), .Y(\U3/U85/Z_26 ) );
  OAI21X1 U3114 ( .A(n3477), .B(n4058), .C(n3476), .Y(\U3/U85/Z_25 ) );
  OAI21X1 U3115 ( .A(n3477), .B(n4056), .C(n3476), .Y(\U3/U85/Z_24 ) );
  OAI21X1 U3116 ( .A(n3477), .B(n4054), .C(n3476), .Y(\U3/U85/Z_23 ) );
  OAI21X1 U3117 ( .A(n3477), .B(n4052), .C(n3476), .Y(\U3/U85/Z_22 ) );
  OAI21X1 U3118 ( .A(n3477), .B(n4050), .C(n3476), .Y(\U3/U85/Z_21 ) );
  OAI21X1 U3119 ( .A(n3477), .B(n4048), .C(n3476), .Y(\U3/U85/Z_20 ) );
  OAI21X1 U3120 ( .A(n3477), .B(n6106), .C(n6107), .Y(\U3/U85/Z_2 ) );
  AOI21X1 U3121 ( .A(\regX[22][2] ), .B(n7253), .C(n3483), .Y(n6107) );
  OAI21X1 U3122 ( .A(n3477), .B(n4046), .C(n3476), .Y(\U3/U85/Z_19 ) );
  OAI21X1 U3123 ( .A(n3477), .B(n4044), .C(n3476), .Y(\U3/U85/Z_18 ) );
  OAI21X1 U3124 ( .A(n3477), .B(n4042), .C(n3476), .Y(\U3/U85/Z_17 ) );
  OAI21X1 U3125 ( .A(n3477), .B(n4040), .C(n3476), .Y(\U3/U85/Z_16 ) );
  OAI21X1 U3126 ( .A(n3477), .B(n4038), .C(n3476), .Y(\U3/U85/Z_15 ) );
  OAI21X1 U3127 ( .A(n3477), .B(n4036), .C(n3476), .Y(\U3/U85/Z_14 ) );
  OAI21X1 U3128 ( .A(n3477), .B(n4034), .C(n3476), .Y(\U3/U85/Z_13 ) );
  OAI21X1 U3129 ( .A(n3477), .B(n4032), .C(n3476), .Y(\U3/U85/Z_12 ) );
  OAI21X1 U3130 ( .A(n3477), .B(n4030), .C(n3476), .Y(\U3/U85/Z_11 ) );
  OAI21X1 U3131 ( .A(n3477), .B(n4028), .C(n3476), .Y(\U3/U85/Z_10 ) );
  OAI21X1 U3132 ( .A(n3477), .B(n6108), .C(n6109), .Y(\U3/U85/Z_1 ) );
  AOI21X1 U3133 ( .A(\regX[22][1] ), .B(n7253), .C(n3483), .Y(n6109) );
  OAI22X1 U3134 ( .A(n3477), .B(n6110), .C(n3475), .D(n3600), .Y(\U3/U85/Z_0 )
         );
  OAI21X1 U3135 ( .A(n3476), .B(n3794), .C(n3477), .Y(\U3/U84/Z_7 ) );
  OAI21X1 U3136 ( .A(n3476), .B(n3793), .C(n3477), .Y(\U3/U84/Z_6 ) );
  OAI21X1 U3137 ( .A(n3476), .B(n3792), .C(n3477), .Y(\U3/U84/Z_5 ) );
  OAI21X1 U3138 ( .A(n3476), .B(n3791), .C(n3477), .Y(\U3/U84/Z_4 ) );
  OAI21X1 U3139 ( .A(n3476), .B(n3790), .C(n3477), .Y(\U3/U84/Z_3 ) );
  INVX1 U3140 ( .A(\regX[11][3] ), .Y(n3790) );
  OAI21X1 U3141 ( .A(n3476), .B(n3789), .C(n3475), .Y(\U3/U84/Z_2 ) );
  INVX1 U3142 ( .A(\regX[11][2] ), .Y(n3789) );
  OAI21X1 U3143 ( .A(n3476), .B(n3788), .C(n3477), .Y(\U3/U84/Z_1 ) );
  INVX1 U3144 ( .A(\regX[11][1] ), .Y(n3788) );
  OAI21X1 U3145 ( .A(n3476), .B(n3786), .C(n3477), .Y(\U3/U84/Z_0 ) );
  INVX1 U3146 ( .A(\regX[11][0] ), .Y(n3786) );
  OAI21X1 U3147 ( .A(n3480), .B(n4026), .C(n6111), .Y(\U3/U82/Z_9 ) );
  AOI22X1 U3148 ( .A(Gy[9]), .B(n7241), .C(N2245), .D(n4257), .Y(n6111) );
  OAI21X1 U3149 ( .A(n3480), .B(n4023), .C(n6112), .Y(\U3/U82/Z_8 ) );
  AOI22X1 U3150 ( .A(Gy[8]), .B(n7241), .C(N2244), .D(n4257), .Y(n6112) );
  OAI21X1 U3151 ( .A(n3480), .B(n6096), .C(n6113), .Y(\U3/U82/Z_7 ) );
  AOI22X1 U3152 ( .A(Gy[7]), .B(n7241), .C(N2243), .D(n4257), .Y(n6113) );
  OAI21X1 U3153 ( .A(n3480), .B(n6098), .C(n6114), .Y(\U3/U82/Z_6 ) );
  AOI22X1 U3154 ( .A(Gy[6]), .B(n7241), .C(N2242), .D(n4257), .Y(n6114) );
  OAI21X1 U3155 ( .A(n5725), .B(n6100), .C(n6115), .Y(\U3/U82/Z_5 ) );
  AOI22X1 U3156 ( .A(Gy[5]), .B(n7241), .C(N2241), .D(n4257), .Y(n6115) );
  OAI21X1 U3157 ( .A(n5725), .B(n6102), .C(n6116), .Y(\U3/U82/Z_4 ) );
  AOI22X1 U3158 ( .A(Gy[4]), .B(n7241), .C(N2240), .D(n4257), .Y(n6116) );
  OAI21X1 U3159 ( .A(n5725), .B(n4070), .C(n6117), .Y(\U3/U82/Z_31 ) );
  AOI21X1 U3160 ( .A(N2267), .B(n4257), .C(n7241), .Y(n6117) );
  OAI21X1 U3161 ( .A(n5725), .B(n4068), .C(n6118), .Y(\U3/U82/Z_30 ) );
  AOI22X1 U3162 ( .A(Gy[30]), .B(n7241), .C(N2266), .D(n4257), .Y(n6118) );
  OAI21X1 U3163 ( .A(n5725), .B(n6104), .C(n6119), .Y(\U3/U82/Z_3 ) );
  AOI22X1 U3164 ( .A(Gy[3]), .B(n7241), .C(N2239), .D(n4257), .Y(n6119) );
  OAI21X1 U3165 ( .A(n5725), .B(n4066), .C(n6120), .Y(\U3/U82/Z_29 ) );
  AOI22X1 U3166 ( .A(Gy[29]), .B(n7241), .C(N2265), .D(n4257), .Y(n6120) );
  OAI21X1 U3167 ( .A(n5725), .B(n4064), .C(n6121), .Y(\U3/U82/Z_28 ) );
  AOI22X1 U3168 ( .A(Gy[28]), .B(n7241), .C(N2264), .D(n4257), .Y(n6121) );
  OAI21X1 U3169 ( .A(n5725), .B(n4062), .C(n6122), .Y(\U3/U82/Z_27 ) );
  AOI22X1 U3170 ( .A(Gy[27]), .B(n7241), .C(N2263), .D(n4257), .Y(n6122) );
  OAI21X1 U3171 ( .A(n5725), .B(n4060), .C(n6123), .Y(\U3/U82/Z_26 ) );
  AOI22X1 U3172 ( .A(Gy[26]), .B(n7241), .C(N2262), .D(n4257), .Y(n6123) );
  OAI21X1 U3173 ( .A(n5725), .B(n4058), .C(n6124), .Y(\U3/U82/Z_25 ) );
  AOI22X1 U3174 ( .A(Gy[25]), .B(n7241), .C(N2261), .D(n4257), .Y(n6124) );
  OAI21X1 U3175 ( .A(n5725), .B(n4056), .C(n6125), .Y(\U3/U82/Z_24 ) );
  AOI22X1 U3176 ( .A(Gy[24]), .B(n7241), .C(N2260), .D(n4257), .Y(n6125) );
  OAI21X1 U3177 ( .A(n5725), .B(n4054), .C(n6126), .Y(\U3/U82/Z_23 ) );
  AOI22X1 U3178 ( .A(Gy[23]), .B(n7241), .C(N2259), .D(n4257), .Y(n6126) );
  OAI21X1 U3179 ( .A(n5725), .B(n4052), .C(n6127), .Y(\U3/U82/Z_22 ) );
  AOI22X1 U3180 ( .A(Gy[22]), .B(n7241), .C(N2258), .D(n4257), .Y(n6127) );
  OAI21X1 U3181 ( .A(n5725), .B(n4050), .C(n6128), .Y(\U3/U82/Z_21 ) );
  AOI22X1 U3182 ( .A(Gy[21]), .B(n7241), .C(N2257), .D(n4257), .Y(n6128) );
  OAI21X1 U3183 ( .A(n5725), .B(n4048), .C(n6129), .Y(\U3/U82/Z_20 ) );
  AOI22X1 U3184 ( .A(Gy[20]), .B(n7241), .C(N2256), .D(n4257), .Y(n6129) );
  OAI21X1 U3185 ( .A(n5725), .B(n6106), .C(n6130), .Y(\U3/U82/Z_2 ) );
  AOI22X1 U3186 ( .A(Gy[2]), .B(n7241), .C(N2238), .D(n4257), .Y(n6130) );
  OAI21X1 U3187 ( .A(n5725), .B(n4046), .C(n6131), .Y(\U3/U82/Z_19 ) );
  AOI22X1 U3188 ( .A(Gy[19]), .B(n7241), .C(N2255), .D(n4257), .Y(n6131) );
  OAI21X1 U3189 ( .A(n5725), .B(n4044), .C(n6132), .Y(\U3/U82/Z_18 ) );
  AOI22X1 U3190 ( .A(Gy[18]), .B(n7241), .C(N2254), .D(n4257), .Y(n6132) );
  OAI21X1 U3191 ( .A(n5725), .B(n4042), .C(n6133), .Y(\U3/U82/Z_17 ) );
  AOI22X1 U3192 ( .A(Gy[17]), .B(n7241), .C(N2253), .D(n4257), .Y(n6133) );
  OAI21X1 U3193 ( .A(n5725), .B(n4040), .C(n6134), .Y(\U3/U82/Z_16 ) );
  AOI22X1 U3194 ( .A(Gy[16]), .B(n7241), .C(N2252), .D(n4257), .Y(n6134) );
  OAI21X1 U3195 ( .A(n5725), .B(n4038), .C(n6135), .Y(\U3/U82/Z_15 ) );
  AOI22X1 U3196 ( .A(Gy[15]), .B(n7241), .C(N2251), .D(n4257), .Y(n6135) );
  OAI21X1 U3197 ( .A(n5725), .B(n4036), .C(n6136), .Y(\U3/U82/Z_14 ) );
  AOI22X1 U3198 ( .A(Gy[14]), .B(n7241), .C(N2250), .D(n4257), .Y(n6136) );
  OAI21X1 U3199 ( .A(n5725), .B(n4034), .C(n6137), .Y(\U3/U82/Z_13 ) );
  AOI22X1 U3200 ( .A(Gy[13]), .B(n7241), .C(N2249), .D(n4257), .Y(n6137) );
  OAI21X1 U3201 ( .A(n5725), .B(n4032), .C(n6138), .Y(\U3/U82/Z_12 ) );
  AOI22X1 U3202 ( .A(Gy[12]), .B(n7241), .C(N2248), .D(n4257), .Y(n6138) );
  OAI21X1 U3203 ( .A(n5725), .B(n4030), .C(n6139), .Y(\U3/U82/Z_11 ) );
  AOI22X1 U3204 ( .A(Gy[11]), .B(n7241), .C(N2247), .D(n4257), .Y(n6139) );
  OAI21X1 U3205 ( .A(n5725), .B(n4028), .C(n6140), .Y(\U3/U82/Z_10 ) );
  AOI22X1 U3206 ( .A(Gy[10]), .B(n7241), .C(N2246), .D(n4257), .Y(n6140) );
  OAI21X1 U3207 ( .A(n5725), .B(n6108), .C(n6141), .Y(\U3/U82/Z_1 ) );
  AOI22X1 U3208 ( .A(Gy[1]), .B(n7241), .C(N2237), .D(n4257), .Y(n6141) );
  OAI21X1 U3209 ( .A(n5725), .B(n6110), .C(n6142), .Y(\U3/U82/Z_0 ) );
  AOI22X1 U3210 ( .A(Gy[0]), .B(n7241), .C(N2236), .D(n4257), .Y(n6142) );
  INVX1 U3211 ( .A(fGx[0]), .Y(n6110) );
  NOR2X1 U3212 ( .A(n3479), .B(n3784), .Y(\U3/U81/Z_7 ) );
  NOR2X1 U3213 ( .A(n3479), .B(n3783), .Y(\U3/U81/Z_6 ) );
  NOR2X1 U3214 ( .A(n3479), .B(n3782), .Y(\U3/U81/Z_5 ) );
  NOR2X1 U3215 ( .A(n3479), .B(n3781), .Y(\U3/U81/Z_4 ) );
  NOR2X1 U3216 ( .A(n3479), .B(n3780), .Y(\U3/U81/Z_3 ) );
  NOR2X1 U3217 ( .A(n3479), .B(n3779), .Y(\U3/U81/Z_2 ) );
  NOR2X1 U3218 ( .A(n3479), .B(n3778), .Y(\U3/U81/Z_1 ) );
  NOR2X1 U3219 ( .A(n3548), .B(n3776), .Y(\U3/U81/Z_0 ) );
  OAI21X1 U3220 ( .A(n3471), .B(n5744), .C(n6143), .Y(\U3/U79/Z_9 ) );
  NAND2X1 U3221 ( .A(N2277), .B(n4257), .Y(n6143) );
  INVX1 U3222 ( .A(Gx[9]), .Y(n5744) );
  OAI21X1 U3223 ( .A(n3471), .B(n5742), .C(n6144), .Y(\U3/U79/Z_8 ) );
  NAND2X1 U3224 ( .A(N2276), .B(n4257), .Y(n6144) );
  INVX1 U3225 ( .A(Gx[8]), .Y(n5742) );
  OAI21X1 U3226 ( .A(n3471), .B(n5740), .C(n6145), .Y(\U3/U79/Z_7 ) );
  NAND2X1 U3227 ( .A(N2275), .B(n4257), .Y(n6145) );
  INVX1 U3228 ( .A(Gx[7]), .Y(n5740) );
  OAI21X1 U3229 ( .A(n3471), .B(n5738), .C(n6146), .Y(\U3/U79/Z_6 ) );
  NAND2X1 U3230 ( .A(N2274), .B(n4257), .Y(n6146) );
  INVX1 U3231 ( .A(Gx[6]), .Y(n5738) );
  OAI21X1 U3232 ( .A(n3471), .B(n5736), .C(n6147), .Y(\U3/U79/Z_5 ) );
  NAND2X1 U3233 ( .A(N2273), .B(n4257), .Y(n6147) );
  INVX1 U3234 ( .A(Gx[5]), .Y(n5736) );
  OAI21X1 U3235 ( .A(n3471), .B(n5734), .C(n6148), .Y(\U3/U79/Z_4 ) );
  NAND2X1 U3236 ( .A(N2272), .B(n4257), .Y(n6148) );
  INVX1 U3237 ( .A(Gx[4]), .Y(n5734) );
  OAI21X1 U3238 ( .A(n3471), .B(n5788), .C(n6149), .Y(\U3/U79/Z_31 ) );
  NAND2X1 U3239 ( .A(N2299), .B(n4257), .Y(n6149) );
  INVX1 U3240 ( .A(Gx[31]), .Y(n5788) );
  OAI21X1 U3241 ( .A(n3471), .B(n5786), .C(n6150), .Y(\U3/U79/Z_30 ) );
  NAND2X1 U3242 ( .A(N2298), .B(n4257), .Y(n6150) );
  INVX1 U3243 ( .A(Gx[30]), .Y(n5786) );
  OAI21X1 U3244 ( .A(n3471), .B(n5732), .C(n6151), .Y(\U3/U79/Z_3 ) );
  NAND2X1 U3245 ( .A(N2271), .B(n4257), .Y(n6151) );
  INVX1 U3246 ( .A(Gx[3]), .Y(n5732) );
  OAI21X1 U3247 ( .A(n3471), .B(n5784), .C(n6152), .Y(\U3/U79/Z_29 ) );
  NAND2X1 U3248 ( .A(N2297), .B(n4257), .Y(n6152) );
  INVX1 U3249 ( .A(Gx[29]), .Y(n5784) );
  OAI21X1 U3250 ( .A(n3471), .B(n5782), .C(n6153), .Y(\U3/U79/Z_28 ) );
  NAND2X1 U3251 ( .A(N2296), .B(n4257), .Y(n6153) );
  INVX1 U3252 ( .A(Gx[28]), .Y(n5782) );
  OAI21X1 U3253 ( .A(n3471), .B(n5780), .C(n6154), .Y(\U3/U79/Z_27 ) );
  NAND2X1 U3254 ( .A(N2295), .B(n4257), .Y(n6154) );
  INVX1 U3255 ( .A(Gx[27]), .Y(n5780) );
  OAI21X1 U3256 ( .A(n3471), .B(n5778), .C(n6155), .Y(\U3/U79/Z_26 ) );
  NAND2X1 U3257 ( .A(N2294), .B(n4257), .Y(n6155) );
  INVX1 U3258 ( .A(Gx[26]), .Y(n5778) );
  OAI21X1 U3259 ( .A(n3471), .B(n5776), .C(n6156), .Y(\U3/U79/Z_25 ) );
  NAND2X1 U3260 ( .A(N2293), .B(n4257), .Y(n6156) );
  INVX1 U3261 ( .A(Gx[25]), .Y(n5776) );
  OAI21X1 U3262 ( .A(n3471), .B(n5774), .C(n6157), .Y(\U3/U79/Z_24 ) );
  NAND2X1 U3263 ( .A(N2292), .B(n4257), .Y(n6157) );
  INVX1 U3264 ( .A(Gx[24]), .Y(n5774) );
  OAI21X1 U3265 ( .A(n3471), .B(n5772), .C(n6158), .Y(\U3/U79/Z_23 ) );
  NAND2X1 U3266 ( .A(N2291), .B(n4257), .Y(n6158) );
  INVX1 U3267 ( .A(Gx[23]), .Y(n5772) );
  OAI21X1 U3268 ( .A(n3471), .B(n5770), .C(n6159), .Y(\U3/U79/Z_22 ) );
  NAND2X1 U3269 ( .A(N2290), .B(n4257), .Y(n6159) );
  INVX1 U3270 ( .A(Gx[22]), .Y(n5770) );
  OAI21X1 U3271 ( .A(n3471), .B(n5768), .C(n6160), .Y(\U3/U79/Z_21 ) );
  NAND2X1 U3272 ( .A(N2289), .B(n4257), .Y(n6160) );
  INVX1 U3273 ( .A(Gx[21]), .Y(n5768) );
  OAI21X1 U3274 ( .A(n3471), .B(n5766), .C(n6161), .Y(\U3/U79/Z_20 ) );
  NAND2X1 U3275 ( .A(N2288), .B(n4257), .Y(n6161) );
  INVX1 U3276 ( .A(Gx[20]), .Y(n5766) );
  OAI21X1 U3277 ( .A(n3471), .B(n5730), .C(n6162), .Y(\U3/U79/Z_2 ) );
  NAND2X1 U3278 ( .A(N2270), .B(n4257), .Y(n6162) );
  INVX1 U3279 ( .A(Gx[2]), .Y(n5730) );
  OAI21X1 U3280 ( .A(n3471), .B(n5764), .C(n6163), .Y(\U3/U79/Z_19 ) );
  NAND2X1 U3281 ( .A(N2287), .B(n4257), .Y(n6163) );
  INVX1 U3282 ( .A(Gx[19]), .Y(n5764) );
  OAI21X1 U3283 ( .A(n3471), .B(n5762), .C(n6164), .Y(\U3/U79/Z_18 ) );
  NAND2X1 U3284 ( .A(N2286), .B(n4257), .Y(n6164) );
  INVX1 U3285 ( .A(Gx[18]), .Y(n5762) );
  OAI21X1 U3286 ( .A(n3471), .B(n5760), .C(n6165), .Y(\U3/U79/Z_17 ) );
  NAND2X1 U3287 ( .A(N2285), .B(n4257), .Y(n6165) );
  INVX1 U3288 ( .A(Gx[17]), .Y(n5760) );
  OAI21X1 U3289 ( .A(n3471), .B(n5758), .C(n6166), .Y(\U3/U79/Z_16 ) );
  NAND2X1 U3290 ( .A(N2284), .B(n4257), .Y(n6166) );
  INVX1 U3291 ( .A(Gx[16]), .Y(n5758) );
  OAI21X1 U3292 ( .A(n3471), .B(n5756), .C(n6167), .Y(\U3/U79/Z_15 ) );
  NAND2X1 U3293 ( .A(N2283), .B(n4257), .Y(n6167) );
  INVX1 U3294 ( .A(Gx[15]), .Y(n5756) );
  OAI21X1 U3295 ( .A(n3471), .B(n5754), .C(n6168), .Y(\U3/U79/Z_14 ) );
  NAND2X1 U3296 ( .A(N2282), .B(n4257), .Y(n6168) );
  INVX1 U3297 ( .A(Gx[14]), .Y(n5754) );
  OAI21X1 U3298 ( .A(n3471), .B(n5752), .C(n6169), .Y(\U3/U79/Z_13 ) );
  NAND2X1 U3299 ( .A(N2281), .B(n4257), .Y(n6169) );
  INVX1 U3300 ( .A(Gx[13]), .Y(n5752) );
  OAI21X1 U3301 ( .A(n3471), .B(n5750), .C(n6170), .Y(\U3/U79/Z_12 ) );
  NAND2X1 U3302 ( .A(N2280), .B(n4257), .Y(n6170) );
  INVX1 U3303 ( .A(Gx[12]), .Y(n5750) );
  OAI21X1 U3304 ( .A(n3471), .B(n5748), .C(n6171), .Y(\U3/U79/Z_11 ) );
  NAND2X1 U3305 ( .A(N2279), .B(n4257), .Y(n6171) );
  INVX1 U3306 ( .A(Gx[11]), .Y(n5748) );
  OAI21X1 U3307 ( .A(n3471), .B(n5746), .C(n6172), .Y(\U3/U79/Z_10 ) );
  NAND2X1 U3308 ( .A(N2278), .B(n4257), .Y(n6172) );
  INVX1 U3309 ( .A(Gx[10]), .Y(n5746) );
  OAI21X1 U3310 ( .A(n3471), .B(n5728), .C(n6173), .Y(\U3/U79/Z_1 ) );
  NAND2X1 U3311 ( .A(N2269), .B(n4257), .Y(n6173) );
  INVX1 U3312 ( .A(Gx[1]), .Y(n5728) );
  OAI21X1 U3313 ( .A(n3471), .B(n5726), .C(n6174), .Y(\U3/U79/Z_0 ) );
  NAND2X1 U3314 ( .A(N2268), .B(n4257), .Y(n6174) );
  INVX1 U3315 ( .A(Gx[0]), .Y(n5726) );
  INVX1 U3316 ( .A(n3547), .Y(n4127) );
  NOR2X1 U3317 ( .A(n3548), .B(n6175), .Y(\U3/U78/Z_9 ) );
  AND2X1 U3318 ( .A(n4257), .B(N2753), .Y(\U3/U78/Z_8 ) );
  AND2X1 U3319 ( .A(n4257), .B(N2752), .Y(\U3/U78/Z_7 ) );
  AND2X1 U3320 ( .A(n4257), .B(N2751), .Y(\U3/U78/Z_6 ) );
  AND2X1 U3321 ( .A(n4257), .B(N2750), .Y(\U3/U78/Z_5 ) );
  NOR2X1 U3322 ( .A(n3548), .B(n6176), .Y(\U3/U78/Z_4 ) );
  NOR2X1 U3323 ( .A(n3548), .B(n6177), .Y(\U3/U78/Z_31 ) );
  NOR2X1 U3324 ( .A(n3548), .B(n6178), .Y(\U3/U78/Z_30 ) );
  NOR2X1 U3325 ( .A(n3548), .B(n6179), .Y(\U3/U78/Z_3 ) );
  NOR2X1 U3326 ( .A(n3548), .B(n6180), .Y(\U3/U78/Z_29 ) );
  NOR2X1 U3327 ( .A(n3548), .B(n6181), .Y(\U3/U78/Z_28 ) );
  NOR2X1 U3328 ( .A(n3548), .B(n6182), .Y(\U3/U78/Z_27 ) );
  NOR2X1 U3329 ( .A(n3548), .B(n6183), .Y(\U3/U78/Z_26 ) );
  NOR2X1 U3330 ( .A(n3548), .B(n6184), .Y(\U3/U78/Z_25 ) );
  NOR2X1 U3331 ( .A(n3548), .B(n6185), .Y(\U3/U78/Z_24 ) );
  NOR2X1 U3332 ( .A(n3548), .B(n6186), .Y(\U3/U78/Z_23 ) );
  NOR2X1 U3333 ( .A(n3548), .B(n6187), .Y(\U3/U78/Z_22 ) );
  NOR2X1 U3334 ( .A(n3548), .B(n6188), .Y(\U3/U78/Z_21 ) );
  NOR2X1 U3335 ( .A(n3548), .B(n6189), .Y(\U3/U78/Z_20 ) );
  NOR2X1 U3336 ( .A(n3548), .B(n6190), .Y(\U3/U78/Z_2 ) );
  NOR2X1 U3337 ( .A(n3548), .B(n6191), .Y(\U3/U78/Z_19 ) );
  NOR2X1 U3338 ( .A(n3548), .B(n6192), .Y(\U3/U78/Z_18 ) );
  NOR2X1 U3339 ( .A(n3548), .B(n6193), .Y(\U3/U78/Z_17 ) );
  NOR2X1 U3340 ( .A(n3548), .B(n6194), .Y(\U3/U78/Z_16 ) );
  NOR2X1 U3341 ( .A(n3548), .B(n6195), .Y(\U3/U78/Z_15 ) );
  NOR2X1 U3342 ( .A(n3548), .B(n6196), .Y(\U3/U78/Z_14 ) );
  NOR2X1 U3343 ( .A(n3548), .B(n6197), .Y(\U3/U78/Z_13 ) );
  NOR2X1 U3344 ( .A(n3548), .B(n6198), .Y(\U3/U78/Z_12 ) );
  NOR2X1 U3345 ( .A(n3548), .B(n6199), .Y(\U3/U78/Z_11 ) );
  NOR2X1 U3346 ( .A(n3548), .B(n6200), .Y(\U3/U78/Z_10 ) );
  NOR2X1 U3347 ( .A(n3548), .B(n6201), .Y(\U3/U78/Z_1 ) );
  AND2X1 U3348 ( .A(n4257), .B(N2648), .Y(\U3/U78/Z_0 ) );
  AND2X1 U3349 ( .A(\U3/U77/DATA2_31 ), .B(n3484), .Y(\U3/U77/Z_31 ) );
  AND2X1 U3350 ( .A(\U3/U77/DATA2_30 ), .B(n3484), .Y(\U3/U77/Z_30 ) );
  AND2X1 U3351 ( .A(\U3/U77/DATA2_29 ), .B(n3484), .Y(\U3/U77/Z_29 ) );
  AND2X1 U3352 ( .A(\U3/U77/DATA2_28 ), .B(n3484), .Y(\U3/U77/Z_28 ) );
  AND2X1 U3353 ( .A(\U3/U77/DATA2_27 ), .B(n3484), .Y(\U3/U77/Z_27 ) );
  AND2X1 U3354 ( .A(\U3/U77/DATA2_26 ), .B(n3484), .Y(\U3/U77/Z_26 ) );
  AND2X1 U3355 ( .A(\U3/U77/DATA2_25 ), .B(n3484), .Y(\U3/U77/Z_25 ) );
  AND2X1 U3356 ( .A(\U3/U77/DATA2_24 ), .B(n3484), .Y(\U3/U77/Z_24 ) );
  AND2X1 U3357 ( .A(\U3/U77/DATA2_23 ), .B(n3484), .Y(\U3/U77/Z_23 ) );
  AND2X1 U3358 ( .A(\U3/U77/DATA2_22 ), .B(n3484), .Y(\U3/U77/Z_22 ) );
  AND2X1 U3359 ( .A(\U3/U77/DATA2_21 ), .B(n3484), .Y(\U3/U77/Z_21 ) );
  AND2X1 U3360 ( .A(\U3/U77/DATA2_20 ), .B(n3484), .Y(\U3/U77/Z_20 ) );
  AND2X1 U3361 ( .A(\U3/U77/DATA2_19 ), .B(n3484), .Y(\U3/U77/Z_19 ) );
  AND2X1 U3362 ( .A(\U3/U77/DATA2_18 ), .B(n3484), .Y(\U3/U77/Z_18 ) );
  AND2X1 U3363 ( .A(\U3/U77/DATA2_17 ), .B(n3484), .Y(\U3/U77/Z_17 ) );
  AND2X1 U3364 ( .A(\U3/U77/DATA2_16 ), .B(n3484), .Y(\U3/U77/Z_16 ) );
  AND2X1 U3365 ( .A(\U3/U77/DATA2_15 ), .B(n3484), .Y(\U3/U77/Z_15 ) );
  AND2X1 U3366 ( .A(N2399), .B(n7253), .Y(\U3/U76/Z_14 ) );
  AND2X1 U3367 ( .A(N2398), .B(n7253), .Y(\U3/U76/Z_13 ) );
  AND2X1 U3368 ( .A(N2397), .B(n7253), .Y(\U3/U76/Z_12 ) );
  AND2X1 U3369 ( .A(N2396), .B(n7253), .Y(\U3/U76/Z_11 ) );
  AND2X1 U3370 ( .A(N2395), .B(n7253), .Y(\U3/U76/Z_10 ) );
  AND2X1 U3371 ( .A(N2117), .B(n7253), .Y(\U3/U75/Z_9 ) );
  AND2X1 U3372 ( .A(N2116), .B(n7253), .Y(\U3/U75/Z_8 ) );
  OAI21X1 U3373 ( .A(n3476), .B(n3911), .C(n6202), .Y(\U3/U75/Z_7 ) );
  NAND2X1 U3374 ( .A(N2115), .B(n7253), .Y(n6202) );
  OAI21X1 U3375 ( .A(n3476), .B(n3910), .C(n6203), .Y(\U3/U75/Z_6 ) );
  NAND2X1 U3376 ( .A(N2114), .B(n7253), .Y(n6203) );
  OAI21X1 U3377 ( .A(n3476), .B(n3909), .C(n6204), .Y(\U3/U75/Z_5 ) );
  NAND2X1 U3378 ( .A(N2113), .B(n7253), .Y(n6204) );
  OAI21X1 U3379 ( .A(n3476), .B(n3908), .C(n6205), .Y(\U3/U75/Z_4 ) );
  NAND2X1 U3380 ( .A(N2112), .B(n7253), .Y(n6205) );
  OAI21X1 U3381 ( .A(n3476), .B(n3907), .C(n6206), .Y(\U3/U75/Z_3 ) );
  NAND2X1 U3382 ( .A(N2111), .B(n7253), .Y(n6206) );
  OAI21X1 U3383 ( .A(n3476), .B(n3906), .C(n6207), .Y(\U3/U75/Z_2 ) );
  NAND2X1 U3384 ( .A(N2110), .B(n7253), .Y(n6207) );
  AND2X1 U3385 ( .A(N2122), .B(n7253), .Y(\U3/U75/Z_14 ) );
  AND2X1 U3386 ( .A(N2121), .B(n7253), .Y(\U3/U75/Z_13 ) );
  AND2X1 U3387 ( .A(N2120), .B(n7253), .Y(\U3/U75/Z_12 ) );
  AND2X1 U3388 ( .A(N2119), .B(n7253), .Y(\U3/U75/Z_11 ) );
  AND2X1 U3389 ( .A(N2118), .B(n7253), .Y(\U3/U75/Z_10 ) );
  OAI21X1 U3390 ( .A(n3476), .B(n3905), .C(n6208), .Y(\U3/U75/Z_1 ) );
  NAND2X1 U3391 ( .A(N2109), .B(n7253), .Y(n6208) );
  OAI21X1 U3392 ( .A(n3476), .B(n3903), .C(n6209), .Y(\U3/U75/Z_0 ) );
  NAND2X1 U3393 ( .A(N2108), .B(n7253), .Y(n6209) );
  AND2X1 U3394 ( .A(n3484), .B(N2267), .Y(\U3/U74/Z_31 ) );
  AND2X1 U3395 ( .A(n3484), .B(N2266), .Y(\U3/U74/Z_30 ) );
  AND2X1 U3396 ( .A(n3484), .B(N2265), .Y(\U3/U74/Z_29 ) );
  AND2X1 U3397 ( .A(n3483), .B(N2264), .Y(\U3/U74/Z_28 ) );
  AND2X1 U3398 ( .A(n3483), .B(N2263), .Y(\U3/U74/Z_27 ) );
  AND2X1 U3399 ( .A(n3483), .B(N2262), .Y(\U3/U74/Z_26 ) );
  AND2X1 U3400 ( .A(n3483), .B(N2261), .Y(\U3/U74/Z_25 ) );
  AND2X1 U3401 ( .A(n3483), .B(N2260), .Y(\U3/U74/Z_24 ) );
  AND2X1 U3402 ( .A(n3483), .B(N2259), .Y(\U3/U74/Z_23 ) );
  AND2X1 U3403 ( .A(n3483), .B(N2258), .Y(\U3/U74/Z_22 ) );
  AND2X1 U3404 ( .A(n3483), .B(N2257), .Y(\U3/U74/Z_21 ) );
  AND2X1 U3405 ( .A(n3483), .B(N2256), .Y(\U3/U74/Z_20 ) );
  AND2X1 U3406 ( .A(n3483), .B(N2255), .Y(\U3/U74/Z_19 ) );
  AND2X1 U3407 ( .A(n3483), .B(N2254), .Y(\U3/U74/Z_18 ) );
  AND2X1 U3408 ( .A(n3483), .B(N2253), .Y(\U3/U74/Z_17 ) );
  AND2X1 U3409 ( .A(n3483), .B(N2252), .Y(\U3/U74/Z_16 ) );
  AND2X1 U3410 ( .A(n3483), .B(N2251), .Y(\U3/U74/Z_15 ) );
  NOR2X1 U3411 ( .A(n3476), .B(n5832), .Y(\U3/U73/Z_31 ) );
  INVX1 U3412 ( .A(N2911), .Y(n5832) );
  NOR2X1 U3413 ( .A(n3476), .B(n5834), .Y(\U3/U73/Z_30 ) );
  INVX1 U3414 ( .A(N2910), .Y(n5834) );
  NOR2X1 U3415 ( .A(n3476), .B(n5835), .Y(\U3/U73/Z_29 ) );
  INVX1 U3416 ( .A(N2909), .Y(n5835) );
  NOR2X1 U3417 ( .A(n3476), .B(n5836), .Y(\U3/U73/Z_28 ) );
  INVX1 U3418 ( .A(N2908), .Y(n5836) );
  NOR2X1 U3419 ( .A(n3476), .B(n5837), .Y(\U3/U73/Z_27 ) );
  INVX1 U3420 ( .A(N2907), .Y(n5837) );
  NOR2X1 U3421 ( .A(n3476), .B(n5838), .Y(\U3/U73/Z_26 ) );
  INVX1 U3422 ( .A(N2906), .Y(n5838) );
  NOR2X1 U3423 ( .A(n3476), .B(n5839), .Y(\U3/U73/Z_25 ) );
  INVX1 U3424 ( .A(N2905), .Y(n5839) );
  NOR2X1 U3425 ( .A(n3476), .B(n5840), .Y(\U3/U73/Z_24 ) );
  INVX1 U3426 ( .A(N2904), .Y(n5840) );
  NOR2X1 U3427 ( .A(n3476), .B(n5841), .Y(\U3/U73/Z_23 ) );
  INVX1 U3428 ( .A(N2903), .Y(n5841) );
  NOR2X1 U3429 ( .A(n3476), .B(n5842), .Y(\U3/U73/Z_22 ) );
  INVX1 U3430 ( .A(N2902), .Y(n5842) );
  NOR2X1 U3431 ( .A(n3476), .B(n5843), .Y(\U3/U73/Z_21 ) );
  INVX1 U3432 ( .A(N2901), .Y(n5843) );
  NOR2X1 U3433 ( .A(n3476), .B(n5845), .Y(\U3/U73/Z_20 ) );
  INVX1 U3434 ( .A(N2900), .Y(n5845) );
  NOR2X1 U3435 ( .A(n3476), .B(n5846), .Y(\U3/U73/Z_19 ) );
  INVX1 U3436 ( .A(N2899), .Y(n5846) );
  NOR2X1 U3437 ( .A(n3476), .B(n5847), .Y(\U3/U73/Z_18 ) );
  INVX1 U3438 ( .A(N2898), .Y(n5847) );
  NOR2X1 U3439 ( .A(n3476), .B(n5848), .Y(\U3/U73/Z_17 ) );
  INVX1 U3440 ( .A(N2897), .Y(n5848) );
  NOR2X1 U3441 ( .A(n3476), .B(n5849), .Y(\U3/U73/Z_16 ) );
  INVX1 U3442 ( .A(N2896), .Y(n5849) );
  NOR2X1 U3443 ( .A(n3476), .B(n5850), .Y(\U3/U73/Z_15 ) );
  INVX1 U3444 ( .A(N2895), .Y(n5850) );
  AND2X1 U3445 ( .A(N2840), .B(n3484), .Y(\U3/U72/Z_31 ) );
  AND2X1 U3446 ( .A(N2839), .B(n3484), .Y(\U3/U72/Z_30 ) );
  AND2X1 U3447 ( .A(N2838), .B(n3484), .Y(\U3/U72/Z_29 ) );
  AND2X1 U3448 ( .A(N2837), .B(n3484), .Y(\U3/U72/Z_28 ) );
  AND2X1 U3449 ( .A(N2836), .B(n3484), .Y(\U3/U72/Z_27 ) );
  AND2X1 U3450 ( .A(N2835), .B(n3484), .Y(\U3/U72/Z_26 ) );
  AND2X1 U3451 ( .A(N2834), .B(n3484), .Y(\U3/U72/Z_25 ) );
  AND2X1 U3452 ( .A(N2833), .B(n3484), .Y(\U3/U72/Z_24 ) );
  AND2X1 U3453 ( .A(N2832), .B(n3484), .Y(\U3/U72/Z_23 ) );
  AND2X1 U3454 ( .A(N2831), .B(n3484), .Y(\U3/U72/Z_22 ) );
  AND2X1 U3455 ( .A(N2830), .B(n3484), .Y(\U3/U72/Z_21 ) );
  AND2X1 U3456 ( .A(N2829), .B(n3484), .Y(\U3/U72/Z_20 ) );
  AND2X1 U3457 ( .A(N2828), .B(n3484), .Y(\U3/U72/Z_19 ) );
  AND2X1 U3458 ( .A(N2827), .B(n3484), .Y(\U3/U72/Z_18 ) );
  AND2X1 U3459 ( .A(N2826), .B(n3484), .Y(\U3/U72/Z_17 ) );
  AND2X1 U3460 ( .A(N2825), .B(n3484), .Y(\U3/U72/Z_16 ) );
  AND2X1 U3461 ( .A(N2824), .B(n3484), .Y(\U3/U72/Z_15 ) );
  AND2X1 U3462 ( .A(N2171), .B(n3484), .Y(\U3/U71/Z_31 ) );
  AND2X1 U3463 ( .A(N2170), .B(n3484), .Y(\U3/U71/Z_30 ) );
  AND2X1 U3464 ( .A(N2169), .B(n3484), .Y(\U3/U71/Z_29 ) );
  AND2X1 U3465 ( .A(N2168), .B(n3484), .Y(\U3/U71/Z_28 ) );
  AND2X1 U3466 ( .A(N2167), .B(n3484), .Y(\U3/U71/Z_27 ) );
  AND2X1 U3467 ( .A(N2166), .B(n3484), .Y(\U3/U71/Z_26 ) );
  AND2X1 U3468 ( .A(N2165), .B(n3484), .Y(\U3/U71/Z_25 ) );
  AND2X1 U3469 ( .A(N2164), .B(n3484), .Y(\U3/U71/Z_24 ) );
  AND2X1 U3470 ( .A(N2163), .B(n3484), .Y(\U3/U71/Z_23 ) );
  AND2X1 U3471 ( .A(N2162), .B(n3484), .Y(\U3/U71/Z_22 ) );
  AND2X1 U3472 ( .A(N2161), .B(n3484), .Y(\U3/U71/Z_21 ) );
  AND2X1 U3473 ( .A(N2160), .B(n3484), .Y(\U3/U71/Z_20 ) );
  AND2X1 U3474 ( .A(N2159), .B(n3484), .Y(\U3/U71/Z_19 ) );
  AND2X1 U3475 ( .A(N2158), .B(n3484), .Y(\U3/U71/Z_18 ) );
  AND2X1 U3476 ( .A(N2157), .B(n3484), .Y(\U3/U71/Z_17 ) );
  AND2X1 U3477 ( .A(N2156), .B(n3484), .Y(\U3/U71/Z_16 ) );
  AND2X1 U3478 ( .A(N2155), .B(n3484), .Y(\U3/U71/Z_15 ) );
  NOR2X1 U3479 ( .A(n3476), .B(n3836), .Y(\U3/U70/Z_8 ) );
  OAI22X1 U3480 ( .A(n3475), .B(n3887), .C(n3476), .D(n3835), .Y(\U3/U70/Z_7 )
         );
  OAI22X1 U3481 ( .A(n3475), .B(n3886), .C(n3476), .D(n3834), .Y(\U3/U70/Z_6 )
         );
  OAI22X1 U3482 ( .A(n3475), .B(n3885), .C(n3476), .D(n3833), .Y(\U3/U70/Z_5 )
         );
  OAI22X1 U3483 ( .A(n3475), .B(n3884), .C(n3476), .D(n3832), .Y(\U3/U70/Z_4 )
         );
  OAI22X1 U3484 ( .A(n3475), .B(n3883), .C(n3476), .D(n3831), .Y(\U3/U70/Z_3 )
         );
  OAI22X1 U3485 ( .A(n3475), .B(n3882), .C(n3476), .D(n3830), .Y(\U3/U70/Z_2 )
         );
  OAI22X1 U3486 ( .A(n3475), .B(n3881), .C(n3476), .D(n3828), .Y(\U3/U70/Z_1 )
         );
  NOR2X1 U3487 ( .A(n3475), .B(n3879), .Y(\U3/U70/Z_0 ) );
  AND2X1 U3488 ( .A(N1352), .B(n7253), .Y(\U3/U69/Z_9 ) );
  AND2X1 U3489 ( .A(N1351), .B(n7253), .Y(\U3/U69/Z_8 ) );
  OAI21X1 U3490 ( .A(n3476), .B(n3911), .C(n6210), .Y(\U3/U69/Z_7 ) );
  NAND2X1 U3491 ( .A(N1350), .B(n7253), .Y(n6210) );
  OAI21X1 U3492 ( .A(n3476), .B(n3910), .C(n6211), .Y(\U3/U69/Z_6 ) );
  NAND2X1 U3493 ( .A(N1349), .B(n7253), .Y(n6211) );
  OAI21X1 U3494 ( .A(n3476), .B(n3909), .C(n6212), .Y(\U3/U69/Z_5 ) );
  NAND2X1 U3495 ( .A(N1348), .B(n7253), .Y(n6212) );
  OAI21X1 U3496 ( .A(n3476), .B(n3908), .C(n6213), .Y(\U3/U69/Z_4 ) );
  NAND2X1 U3497 ( .A(N1347), .B(n7253), .Y(n6213) );
  OAI21X1 U3498 ( .A(n3476), .B(n3907), .C(n6214), .Y(\U3/U69/Z_3 ) );
  NAND2X1 U3499 ( .A(N1346), .B(n7253), .Y(n6214) );
  OAI21X1 U3500 ( .A(n3476), .B(n3906), .C(n6215), .Y(\U3/U69/Z_2 ) );
  NAND2X1 U3501 ( .A(N1345), .B(n7253), .Y(n6215) );
  AND2X1 U3502 ( .A(N1356), .B(n7253), .Y(\U3/U69/Z_13 ) );
  AND2X1 U3503 ( .A(N1355), .B(n7253), .Y(\U3/U69/Z_12 ) );
  AND2X1 U3504 ( .A(N1354), .B(n7253), .Y(\U3/U69/Z_11 ) );
  AND2X1 U3505 ( .A(N1353), .B(n7253), .Y(\U3/U69/Z_10 ) );
  OAI21X1 U3506 ( .A(n3476), .B(n3905), .C(n6216), .Y(\U3/U69/Z_1 ) );
  NAND2X1 U3507 ( .A(N1344), .B(n7253), .Y(n6216) );
  OAI21X1 U3508 ( .A(n3476), .B(n3903), .C(n6217), .Y(\U3/U69/Z_0 ) );
  NAND2X1 U3509 ( .A(N1343), .B(n7253), .Y(n6217) );
  AND2X1 U3510 ( .A(N2107), .B(n3484), .Y(\U3/U68/Z_31 ) );
  AND2X1 U3511 ( .A(N2106), .B(n3484), .Y(\U3/U68/Z_30 ) );
  AND2X1 U3512 ( .A(N2105), .B(n3484), .Y(\U3/U68/Z_29 ) );
  AND2X1 U3513 ( .A(N2104), .B(n3484), .Y(\U3/U68/Z_28 ) );
  AND2X1 U3514 ( .A(N2103), .B(n3484), .Y(\U3/U68/Z_27 ) );
  AND2X1 U3515 ( .A(N2102), .B(n3484), .Y(\U3/U68/Z_26 ) );
  AND2X1 U3516 ( .A(N2101), .B(n3484), .Y(\U3/U68/Z_25 ) );
  AND2X1 U3517 ( .A(N2100), .B(n3484), .Y(\U3/U68/Z_24 ) );
  AND2X1 U3518 ( .A(N2099), .B(n3484), .Y(\U3/U68/Z_23 ) );
  AND2X1 U3519 ( .A(N2098), .B(n3484), .Y(\U3/U68/Z_22 ) );
  AND2X1 U3520 ( .A(N2097), .B(n3484), .Y(\U3/U68/Z_21 ) );
  AND2X1 U3521 ( .A(N2096), .B(n3484), .Y(\U3/U68/Z_20 ) );
  AND2X1 U3522 ( .A(N2095), .B(n3484), .Y(\U3/U68/Z_19 ) );
  AND2X1 U3523 ( .A(N2094), .B(n3484), .Y(\U3/U68/Z_18 ) );
  AND2X1 U3524 ( .A(N2093), .B(n3484), .Y(\U3/U68/Z_17 ) );
  AND2X1 U3525 ( .A(N2092), .B(n3484), .Y(\U3/U68/Z_16 ) );
  AND2X1 U3526 ( .A(N2091), .B(n3484), .Y(\U3/U68/Z_15 ) );
  OAI21X1 U3527 ( .A(n3475), .B(n3575), .C(n3476), .Y(\U3/U65/Z_7 ) );
  OAI21X1 U3528 ( .A(n3475), .B(n3573), .C(n3476), .Y(\U3/U65/Z_6 ) );
  OAI21X1 U3529 ( .A(n3475), .B(n3571), .C(n3476), .Y(\U3/U65/Z_5 ) );
  OAI21X1 U3530 ( .A(n3475), .B(n3569), .C(n3476), .Y(\U3/U65/Z_4 ) );
  OAI21X1 U3531 ( .A(n3475), .B(n3567), .C(n3476), .Y(\U3/U65/Z_3 ) );
  OAI21X1 U3532 ( .A(n3475), .B(n3565), .C(n3476), .Y(\U3/U65/Z_2 ) );
  OAI21X1 U3533 ( .A(n3475), .B(n3563), .C(n3476), .Y(\U3/U65/Z_1 ) );
  OAI21X1 U3534 ( .A(n3475), .B(n3560), .C(n3476), .Y(\U3/U65/Z_0 ) );
  NOR2X1 U3535 ( .A(n3476), .B(n3803), .Y(\U3/U64/Z_7 ) );
  NOR2X1 U3536 ( .A(n3476), .B(n3802), .Y(\U3/U64/Z_6 ) );
  NOR2X1 U3537 ( .A(n3476), .B(n3801), .Y(\U3/U64/Z_5 ) );
  NOR2X1 U3538 ( .A(n3476), .B(n3800), .Y(\U3/U64/Z_4 ) );
  NOR2X1 U3539 ( .A(n3476), .B(n3799), .Y(\U3/U64/Z_3 ) );
  NOR2X1 U3540 ( .A(n3476), .B(n3798), .Y(\U3/U64/Z_2 ) );
  NOR2X1 U3541 ( .A(n3476), .B(n3797), .Y(\U3/U64/Z_1 ) );
  OAI21X1 U3542 ( .A(n3476), .B(n3795), .C(n3475), .Y(\U3/U64/Z_0 ) );
  INVX1 U3543 ( .A(N1615), .Y(n3795) );
  NAND2X1 U3544 ( .A(n4257), .B(n4131), .Y(n5791) );
  NOR2X1 U3545 ( .A(n5692), .B(n3640), .Y(\U3/U63/Z_7 ) );
  NOR2X1 U3546 ( .A(n5692), .B(n3639), .Y(\U3/U63/Z_6 ) );
  NOR2X1 U3547 ( .A(n5692), .B(n3638), .Y(\U3/U63/Z_5 ) );
  NOR2X1 U3548 ( .A(n5692), .B(n3637), .Y(\U3/U63/Z_4 ) );
  NOR2X1 U3549 ( .A(n5692), .B(n3636), .Y(\U3/U63/Z_3 ) );
  NAND2X1 U3550 ( .A(bCE), .B(n3635), .Y(\U3/U63/Z_2 ) );
  NOR2X1 U3551 ( .A(n5692), .B(n3634), .Y(\U3/U63/Z_1 ) );
  NAND2X1 U3552 ( .A(bCE), .B(n3632), .Y(\U3/U63/Z_0 ) );
  NAND2X1 U3553 ( .A(N2549), .B(n4080), .Y(\U3/U136/Z_0 ) );
  NOR2X1 U3554 ( .A(n4272), .B(n3966), .Y(\U3/U134/Z_9 ) );
  INVX1 U3555 ( .A(Gy[9]), .Y(n3966) );
  NOR2X1 U3556 ( .A(n4272), .B(n3964), .Y(\U3/U134/Z_8 ) );
  INVX1 U3557 ( .A(Gy[8]), .Y(n3964) );
  NOR2X1 U3558 ( .A(n4272), .B(n3962), .Y(\U3/U134/Z_7 ) );
  INVX1 U3559 ( .A(Gy[7]), .Y(n3962) );
  NOR2X1 U3560 ( .A(n4272), .B(n3960), .Y(\U3/U134/Z_6 ) );
  INVX1 U3561 ( .A(Gy[6]), .Y(n3960) );
  NOR2X1 U3562 ( .A(n4272), .B(n3958), .Y(\U3/U134/Z_5 ) );
  INVX1 U3563 ( .A(Gy[5]), .Y(n3958) );
  NOR2X1 U3564 ( .A(n4272), .B(n3956), .Y(\U3/U134/Z_4 ) );
  INVX1 U3565 ( .A(Gy[4]), .Y(n3956) );
  NOR2X1 U3566 ( .A(n4272), .B(n3954), .Y(\U3/U134/Z_3 ) );
  INVX1 U3567 ( .A(Gy[3]), .Y(n3954) );
  NOR2X1 U3568 ( .A(n4272), .B(n3952), .Y(\U3/U134/Z_2 ) );
  INVX1 U3569 ( .A(Gy[2]), .Y(n3952) );
  NOR2X1 U3570 ( .A(n4272), .B(n3968), .Y(\U3/U134/Z_10 ) );
  INVX1 U3571 ( .A(Gy[10]), .Y(n3968) );
  NOR2X1 U3572 ( .A(n4272), .B(n3950), .Y(\U3/U134/Z_1 ) );
  INVX1 U3573 ( .A(Gy[1]), .Y(n3950) );
  NOR2X1 U3574 ( .A(n4272), .B(n3947), .Y(\U3/U134/Z_0 ) );
  INVX1 U3575 ( .A(Gy[0]), .Y(n3947) );
  INVX1 U3576 ( .A(n3707), .Y(n4272) );
  NAND2X1 U3577 ( .A(n3864), .B(n4128), .Y(n3707) );
  OAI21X1 U3578 ( .A(n3475), .B(n3899), .C(n6218), .Y(\U3/U125/Z_7 ) );
  OAI21X1 U3579 ( .A(n3475), .B(n3898), .C(n6218), .Y(\U3/U125/Z_6 ) );
  OAI21X1 U3580 ( .A(n3475), .B(n3897), .C(n6218), .Y(\U3/U125/Z_5 ) );
  OAI21X1 U3581 ( .A(n3475), .B(n3896), .C(n6218), .Y(\U3/U125/Z_4 ) );
  OAI21X1 U3582 ( .A(n3475), .B(n3895), .C(n6218), .Y(\U3/U125/Z_3 ) );
  OAI21X1 U3583 ( .A(n3475), .B(n3894), .C(n6218), .Y(\U3/U125/Z_2 ) );
  OAI21X1 U3584 ( .A(n3475), .B(n3893), .C(n6218), .Y(\U3/U125/Z_1 ) );
  NAND2X1 U3585 ( .A(dy[1]), .B(n7202), .Y(n6218) );
  OAI22X1 U3586 ( .A(n5161), .B(n5825), .C(n3475), .D(n3891), .Y(\U3/U125/Z_0 ) );
  NAND2X1 U3587 ( .A(n5161), .B(n3475), .Y(\U3/U124/Z_0 ) );
  NOR2X1 U3588 ( .A(n4028), .B(n3482), .Y(\U3/U122/Z_9 ) );
  INVX1 U3589 ( .A(fGx[10]), .Y(n4028) );
  NOR2X1 U3590 ( .A(n4026), .B(n3482), .Y(\U3/U122/Z_8 ) );
  INVX1 U3591 ( .A(fGx[9]), .Y(n4026) );
  OAI21X1 U3592 ( .A(n5826), .B(n4023), .C(n6219), .Y(\U3/U122/Z_7 ) );
  OAI21X1 U3593 ( .A(n6220), .B(n6221), .C(n7205), .Y(n6219) );
  NAND2X1 U3594 ( .A(n6222), .B(n6223), .Y(n6221) );
  NOR2X1 U3595 ( .A(n6224), .B(n6225), .Y(n6223) );
  OAI21X1 U3596 ( .A(n3932), .B(n6226), .C(n6227), .Y(n6225) );
  AOI22X1 U3597 ( .A(n6228), .B(N1382), .C(n6229), .D(N1440), .Y(n6227) );
  OAI21X1 U3598 ( .A(n3875), .B(n6230), .C(n6231), .Y(n6224) );
  AOI22X1 U3599 ( .A(n6232), .B(\regX[3][7] ), .C(n6233), .D(\regX[13][7] ), 
        .Y(n6231) );
  INVX1 U3600 ( .A(\regX[5][7] ), .Y(n3875) );
  NOR2X1 U3601 ( .A(n6234), .B(n6235), .Y(n6222) );
  OAI21X1 U3602 ( .A(n3813), .B(n6236), .C(n6237), .Y(n6235) );
  AOI22X1 U3603 ( .A(n6238), .B(\regX[1][7] ), .C(n6239), .D(\regX[11][7] ), 
        .Y(n6237) );
  OAI21X1 U3604 ( .A(n3836), .B(n6240), .C(n6241), .Y(n6234) );
  AOI22X1 U3605 ( .A(n6242), .B(\regX[8][7] ), .C(n6243), .D(N1622), .Y(n6241)
         );
  NAND2X1 U3606 ( .A(n6244), .B(n6245), .Y(n6220) );
  NOR2X1 U3607 ( .A(n6246), .B(n6247), .Y(n6245) );
  OAI21X1 U3608 ( .A(n3784), .B(n6248), .C(n6249), .Y(n6247) );
  AOI22X1 U3609 ( .A(n6250), .B(\regX[16][7] ), .C(n6251), .D(N1742), .Y(n6249) );
  OAI21X1 U3610 ( .A(n3661), .B(n6252), .C(n6253), .Y(n6246) );
  AOI22X1 U3611 ( .A(n6254), .B(\regX[22][7] ), .C(n6255), .D(\regX[15][7] ), 
        .Y(n6253) );
  NOR2X1 U3612 ( .A(n6256), .B(n6257), .Y(n6244) );
  OAI21X1 U3613 ( .A(n3595), .B(n6258), .C(n6259), .Y(n6257) );
  AOI22X1 U3614 ( .A(n6260), .B(\regX[24][7] ), .C(n6261), .D(\regX[21][7] ), 
        .Y(n6259) );
  OAI21X1 U3615 ( .A(n3640), .B(n6262), .C(n6263), .Y(n6256) );
  AOI22X1 U3616 ( .A(n6264), .B(\regX[20][7] ), .C(n6265), .D(\regX[18][7] ), 
        .Y(n6263) );
  INVX1 U3617 ( .A(\regX[19][7] ), .Y(n3640) );
  INVX1 U3618 ( .A(fGx[8]), .Y(n4023) );
  OAI21X1 U3619 ( .A(n5826), .B(n6096), .C(n6266), .Y(\U3/U122/Z_6 ) );
  OAI21X1 U3620 ( .A(n6267), .B(n6268), .C(n7205), .Y(n6266) );
  NAND2X1 U3621 ( .A(n6269), .B(n6270), .Y(n6268) );
  NOR2X1 U3622 ( .A(n6271), .B(n6272), .Y(n6270) );
  OAI21X1 U3623 ( .A(n3931), .B(n6226), .C(n6273), .Y(n6272) );
  AOI22X1 U3624 ( .A(n6228), .B(N1381), .C(n6229), .D(N1439), .Y(n6273) );
  OAI21X1 U3625 ( .A(n3874), .B(n6230), .C(n6274), .Y(n6271) );
  AOI22X1 U3626 ( .A(n6232), .B(\regX[3][6] ), .C(n6233), .D(\regX[13][6] ), 
        .Y(n6274) );
  INVX1 U3627 ( .A(\regX[5][6] ), .Y(n3874) );
  NOR2X1 U3628 ( .A(n6275), .B(n6276), .Y(n6269) );
  OAI21X1 U3629 ( .A(n3812), .B(n6236), .C(n6277), .Y(n6276) );
  AOI22X1 U3630 ( .A(n6238), .B(\regX[1][6] ), .C(n6239), .D(\regX[11][6] ), 
        .Y(n6277) );
  OAI21X1 U3631 ( .A(n3835), .B(n6240), .C(n6278), .Y(n6275) );
  AOI22X1 U3632 ( .A(n6242), .B(\regX[8][6] ), .C(n6243), .D(N1621), .Y(n6278)
         );
  NAND2X1 U3633 ( .A(n6279), .B(n6280), .Y(n6267) );
  NOR2X1 U3634 ( .A(n6281), .B(n6282), .Y(n6280) );
  OAI21X1 U3635 ( .A(n3783), .B(n6248), .C(n6283), .Y(n6282) );
  AOI22X1 U3636 ( .A(n6250), .B(\regX[16][6] ), .C(n6251), .D(N1741), .Y(n6283) );
  OAI21X1 U3637 ( .A(n3660), .B(n6252), .C(n6284), .Y(n6281) );
  AOI22X1 U3638 ( .A(n6254), .B(\regX[22][6] ), .C(n6255), .D(\regX[15][6] ), 
        .Y(n6284) );
  NOR2X1 U3639 ( .A(n6285), .B(n6286), .Y(n6279) );
  OAI21X1 U3640 ( .A(n3594), .B(n6258), .C(n6287), .Y(n6286) );
  AOI22X1 U3641 ( .A(n6260), .B(\regX[24][6] ), .C(n6261), .D(\regX[21][6] ), 
        .Y(n6287) );
  OAI21X1 U3642 ( .A(n3639), .B(n6262), .C(n6288), .Y(n6285) );
  AOI22X1 U3643 ( .A(n6264), .B(\regX[20][6] ), .C(n6265), .D(\regX[18][6] ), 
        .Y(n6288) );
  INVX1 U3644 ( .A(\regX[19][6] ), .Y(n3639) );
  INVX1 U3645 ( .A(fGx[7]), .Y(n6096) );
  OAI21X1 U3646 ( .A(n5826), .B(n6098), .C(n6289), .Y(\U3/U122/Z_5 ) );
  OAI21X1 U3647 ( .A(n6290), .B(n6291), .C(n7205), .Y(n6289) );
  NAND2X1 U3648 ( .A(n6292), .B(n6293), .Y(n6291) );
  NOR2X1 U3649 ( .A(n6294), .B(n6295), .Y(n6293) );
  OAI21X1 U3650 ( .A(n3930), .B(n6226), .C(n6296), .Y(n6295) );
  AOI22X1 U3651 ( .A(n6228), .B(N1380), .C(n6229), .D(N1438), .Y(n6296) );
  OAI21X1 U3652 ( .A(n3873), .B(n6230), .C(n6297), .Y(n6294) );
  AOI22X1 U3653 ( .A(n6232), .B(\regX[3][5] ), .C(n6233), .D(\regX[13][5] ), 
        .Y(n6297) );
  INVX1 U3654 ( .A(\regX[5][5] ), .Y(n3873) );
  NOR2X1 U3655 ( .A(n6298), .B(n6299), .Y(n6292) );
  OAI21X1 U3656 ( .A(n3811), .B(n6236), .C(n6300), .Y(n6299) );
  AOI22X1 U3657 ( .A(n6238), .B(\regX[1][5] ), .C(n6239), .D(\regX[11][5] ), 
        .Y(n6300) );
  OAI21X1 U3658 ( .A(n3834), .B(n6240), .C(n6301), .Y(n6298) );
  AOI22X1 U3659 ( .A(n6242), .B(\regX[8][5] ), .C(n6243), .D(N1620), .Y(n6301)
         );
  NAND2X1 U3660 ( .A(n6302), .B(n6303), .Y(n6290) );
  NOR2X1 U3661 ( .A(n6304), .B(n6305), .Y(n6303) );
  OAI21X1 U3662 ( .A(n3782), .B(n6248), .C(n6306), .Y(n6305) );
  AOI22X1 U3663 ( .A(n6250), .B(\regX[16][5] ), .C(n6251), .D(N1740), .Y(n6306) );
  OAI21X1 U3664 ( .A(n3659), .B(n6252), .C(n6307), .Y(n6304) );
  AOI22X1 U3665 ( .A(n6254), .B(\regX[22][5] ), .C(n6255), .D(\regX[15][5] ), 
        .Y(n6307) );
  NOR2X1 U3666 ( .A(n6308), .B(n6309), .Y(n6302) );
  OAI21X1 U3667 ( .A(n3593), .B(n6258), .C(n6310), .Y(n6309) );
  AOI22X1 U3668 ( .A(n6260), .B(\regX[24][5] ), .C(n6261), .D(\regX[21][5] ), 
        .Y(n6310) );
  OAI21X1 U3669 ( .A(n3638), .B(n6262), .C(n6311), .Y(n6308) );
  AOI22X1 U3670 ( .A(n6264), .B(\regX[20][5] ), .C(n6265), .D(\regX[18][5] ), 
        .Y(n6311) );
  INVX1 U3671 ( .A(\regX[19][5] ), .Y(n3638) );
  INVX1 U3672 ( .A(fGx[6]), .Y(n6098) );
  OAI21X1 U3673 ( .A(n5826), .B(n6100), .C(n6312), .Y(\U3/U122/Z_4 ) );
  OAI21X1 U3674 ( .A(n6313), .B(n6314), .C(n7205), .Y(n6312) );
  NAND2X1 U3675 ( .A(n6315), .B(n6316), .Y(n6314) );
  NOR2X1 U3676 ( .A(n6317), .B(n6318), .Y(n6316) );
  OAI21X1 U3677 ( .A(n3929), .B(n6226), .C(n6319), .Y(n6318) );
  AOI22X1 U3678 ( .A(n6228), .B(N1379), .C(n6229), .D(N1437), .Y(n6319) );
  INVX1 U3679 ( .A(n6320), .Y(n6229) );
  OAI21X1 U3680 ( .A(n3872), .B(n6230), .C(n6321), .Y(n6317) );
  AOI22X1 U3681 ( .A(n6232), .B(\regX[3][4] ), .C(n6233), .D(\regX[13][4] ), 
        .Y(n6321) );
  INVX1 U3682 ( .A(n6322), .Y(n6232) );
  INVX1 U3683 ( .A(\regX[5][4] ), .Y(n3872) );
  NOR2X1 U3684 ( .A(n6323), .B(n6324), .Y(n6315) );
  OAI21X1 U3685 ( .A(n3810), .B(n6236), .C(n6325), .Y(n6324) );
  AOI22X1 U3686 ( .A(n6238), .B(\regX[1][4] ), .C(n6239), .D(\regX[11][4] ), 
        .Y(n6325) );
  OAI21X1 U3687 ( .A(n3833), .B(n6240), .C(n6326), .Y(n6323) );
  AOI22X1 U3688 ( .A(n6242), .B(\regX[8][4] ), .C(n6243), .D(N1619), .Y(n6326)
         );
  NAND2X1 U3689 ( .A(n6327), .B(n6328), .Y(n6313) );
  NOR2X1 U3690 ( .A(n6329), .B(n6330), .Y(n6328) );
  OAI21X1 U3691 ( .A(n3781), .B(n6248), .C(n6331), .Y(n6330) );
  AOI22X1 U3692 ( .A(n6250), .B(\regX[16][4] ), .C(n6251), .D(N1739), .Y(n6331) );
  OAI21X1 U3693 ( .A(n3658), .B(n6252), .C(n6332), .Y(n6329) );
  AOI22X1 U3694 ( .A(n6254), .B(\regX[22][4] ), .C(n6255), .D(\regX[15][4] ), 
        .Y(n6332) );
  INVX1 U3695 ( .A(n6333), .Y(n6254) );
  NOR2X1 U3696 ( .A(n6334), .B(n6335), .Y(n6327) );
  OAI21X1 U3697 ( .A(n3592), .B(n6258), .C(n6336), .Y(n6335) );
  AOI22X1 U3698 ( .A(n6260), .B(\regX[24][4] ), .C(n6261), .D(\regX[21][4] ), 
        .Y(n6336) );
  INVX1 U3699 ( .A(n6337), .Y(n6261) );
  OAI21X1 U3700 ( .A(n3637), .B(n6262), .C(n6338), .Y(n6334) );
  AOI22X1 U3701 ( .A(n6264), .B(\regX[20][4] ), .C(n6265), .D(\regX[18][4] ), 
        .Y(n6338) );
  INVX1 U3702 ( .A(n6339), .Y(n6264) );
  INVX1 U3703 ( .A(\regX[19][4] ), .Y(n3637) );
  INVX1 U3704 ( .A(fGx[5]), .Y(n6100) );
  OAI21X1 U3705 ( .A(n5826), .B(n6102), .C(n6340), .Y(\U3/U122/Z_3 ) );
  OAI21X1 U3706 ( .A(n6341), .B(n6342), .C(n7205), .Y(n6340) );
  NAND2X1 U3707 ( .A(n6343), .B(n6344), .Y(n6342) );
  NOR2X1 U3708 ( .A(n6345), .B(n6346), .Y(n6344) );
  OAI21X1 U3709 ( .A(n3832), .B(n6240), .C(n6347), .Y(n6346) );
  AOI22X1 U3710 ( .A(n6238), .B(\regX[1][3] ), .C(n6239), .D(\regX[11][3] ), 
        .Y(n6347) );
  INVX1 U3711 ( .A(\regX[7][3] ), .Y(n3832) );
  OAI21X1 U3712 ( .A(n3591), .B(n6258), .C(n6348), .Y(n6345) );
  AOI22X1 U3713 ( .A(n6242), .B(\regX[8][3] ), .C(n6243), .D(N1618), .Y(n6348)
         );
  INVX1 U3714 ( .A(\regX[23][3] ), .Y(n3591) );
  NOR2X1 U3715 ( .A(n6349), .B(n6350), .Y(n6343) );
  OAI21X1 U3716 ( .A(n3809), .B(n6236), .C(n6351), .Y(n6350) );
  AOI22X1 U3717 ( .A(n6352), .B(\regX[5][3] ), .C(n6353), .D(\regX[0][3] ), 
        .Y(n6351) );
  OAI21X1 U3718 ( .A(n3883), .B(n6320), .C(n6354), .Y(n6349) );
  AOI22X1 U3719 ( .A(n6228), .B(N1378), .C(n6233), .D(\regX[13][3] ), .Y(n6354) );
  INVX1 U3720 ( .A(N1436), .Y(n3883) );
  NAND3X1 U3721 ( .A(n6355), .B(n6356), .C(n6357), .Y(n6341) );
  NOR2X1 U3722 ( .A(n6358), .B(n6359), .Y(n6357) );
  OAI21X1 U3723 ( .A(n3657), .B(n6252), .C(n6360), .Y(n6359) );
  AOI22X1 U3724 ( .A(n6255), .B(\regX[15][3] ), .C(n6361), .D(N1680), .Y(n6360) );
  INVX1 U3725 ( .A(\regX[17][3] ), .Y(n3657) );
  OAI21X1 U3726 ( .A(n3636), .B(n6262), .C(n6362), .Y(n6358) );
  AOI22X1 U3727 ( .A(n6250), .B(\regX[16][3] ), .C(n6251), .D(N1738), .Y(n6362) );
  INVX1 U3728 ( .A(\regX[19][3] ), .Y(n3636) );
  NOR2X1 U3729 ( .A(n6363), .B(n6364), .Y(n6356) );
  OAI22X1 U3730 ( .A(n3604), .B(n6333), .C(n3626), .D(n6339), .Y(n6364) );
  INVX1 U3731 ( .A(\regX[20][3] ), .Y(n3626) );
  INVX1 U3732 ( .A(\regX[22][3] ), .Y(n3604) );
  OAI22X1 U3733 ( .A(n3567), .B(n6365), .C(n3845), .D(n6366), .Y(n6363) );
  INVX1 U3734 ( .A(\regX[24][3] ), .Y(n3567) );
  AOI21X1 U3735 ( .A(n6265), .B(\regX[18][3] ), .C(n6367), .Y(n6355) );
  OAI22X1 U3736 ( .A(n3615), .B(n6337), .C(n3895), .D(n6322), .Y(n6367) );
  INVX1 U3737 ( .A(\regX[3][3] ), .Y(n3895) );
  INVX1 U3738 ( .A(fGx[4]), .Y(n6102) );
  NOR2X1 U3739 ( .A(n4068), .B(n3482), .Y(\U3/U122/Z_29 ) );
  INVX1 U3740 ( .A(fGx[30]), .Y(n4068) );
  NOR2X1 U3741 ( .A(n4066), .B(n3482), .Y(\U3/U122/Z_28 ) );
  INVX1 U3742 ( .A(fGx[29]), .Y(n4066) );
  NOR2X1 U3743 ( .A(n4064), .B(n3482), .Y(\U3/U122/Z_27 ) );
  INVX1 U3744 ( .A(fGx[28]), .Y(n4064) );
  NOR2X1 U3745 ( .A(n4062), .B(n3482), .Y(\U3/U122/Z_26 ) );
  INVX1 U3746 ( .A(fGx[27]), .Y(n4062) );
  NOR2X1 U3747 ( .A(n4060), .B(n3482), .Y(\U3/U122/Z_25 ) );
  INVX1 U3748 ( .A(fGx[26]), .Y(n4060) );
  NOR2X1 U3749 ( .A(n4058), .B(n5826), .Y(\U3/U122/Z_24 ) );
  INVX1 U3750 ( .A(fGx[25]), .Y(n4058) );
  NOR2X1 U3751 ( .A(n4056), .B(n5826), .Y(\U3/U122/Z_23 ) );
  INVX1 U3752 ( .A(fGx[24]), .Y(n4056) );
  NOR2X1 U3753 ( .A(n4054), .B(n5826), .Y(\U3/U122/Z_22 ) );
  INVX1 U3754 ( .A(fGx[23]), .Y(n4054) );
  NOR2X1 U3755 ( .A(n4052), .B(n5826), .Y(\U3/U122/Z_21 ) );
  INVX1 U3756 ( .A(fGx[22]), .Y(n4052) );
  NOR2X1 U3757 ( .A(n4050), .B(n5826), .Y(\U3/U122/Z_20 ) );
  INVX1 U3758 ( .A(fGx[21]), .Y(n4050) );
  OAI21X1 U3759 ( .A(n5826), .B(n6104), .C(n6368), .Y(\U3/U122/Z_2 ) );
  OAI21X1 U3760 ( .A(n6369), .B(n6370), .C(n7205), .Y(n6368) );
  NAND2X1 U3761 ( .A(n6371), .B(n6372), .Y(n6370) );
  NOR2X1 U3762 ( .A(n6373), .B(n6374), .Y(n6372) );
  OAI21X1 U3763 ( .A(n3831), .B(n6240), .C(n6375), .Y(n6374) );
  AOI22X1 U3764 ( .A(n6238), .B(\regX[1][2] ), .C(n6239), .D(\regX[11][2] ), 
        .Y(n6375) );
  INVX1 U3765 ( .A(\regX[7][2] ), .Y(n3831) );
  OAI21X1 U3766 ( .A(n3590), .B(n6258), .C(n6376), .Y(n6373) );
  AOI22X1 U3767 ( .A(n6242), .B(\regX[8][2] ), .C(n6243), .D(N1617), .Y(n6376)
         );
  INVX1 U3768 ( .A(\regX[23][2] ), .Y(n3590) );
  NOR2X1 U3769 ( .A(n6377), .B(n6378), .Y(n6371) );
  OAI21X1 U3770 ( .A(n3808), .B(n6236), .C(n6379), .Y(n6378) );
  AOI22X1 U3771 ( .A(n6352), .B(\regX[5][2] ), .C(n6353), .D(\regX[0][2] ), 
        .Y(n6379) );
  OAI21X1 U3772 ( .A(n3882), .B(n6320), .C(n6380), .Y(n6377) );
  AOI22X1 U3773 ( .A(n6228), .B(N1377), .C(n6233), .D(\regX[13][2] ), .Y(n6380) );
  INVX1 U3774 ( .A(N1435), .Y(n3882) );
  NAND3X1 U3775 ( .A(n6381), .B(n6382), .C(n6383), .Y(n6369) );
  NOR2X1 U3776 ( .A(n6384), .B(n6385), .Y(n6383) );
  OAI21X1 U3777 ( .A(n3656), .B(n6252), .C(n6386), .Y(n6385) );
  AOI22X1 U3778 ( .A(n6255), .B(\regX[15][2] ), .C(n6361), .D(N1679), .Y(n6386) );
  INVX1 U3779 ( .A(\regX[17][2] ), .Y(n3656) );
  OAI21X1 U3780 ( .A(n3635), .B(n6262), .C(n6387), .Y(n6384) );
  AOI22X1 U3781 ( .A(n6250), .B(\regX[16][2] ), .C(n6251), .D(N1737), .Y(n6387) );
  INVX1 U3782 ( .A(\regX[19][2] ), .Y(n3635) );
  NOR2X1 U3783 ( .A(n6388), .B(n6389), .Y(n6382) );
  OAI22X1 U3784 ( .A(n3603), .B(n6333), .C(n3625), .D(n6339), .Y(n6389) );
  OAI22X1 U3785 ( .A(n3565), .B(n6365), .C(n3844), .D(n6366), .Y(n6388) );
  AOI21X1 U3786 ( .A(n6265), .B(\regX[18][2] ), .C(n6390), .Y(n6381) );
  OAI22X1 U3787 ( .A(n3614), .B(n6337), .C(n3894), .D(n6322), .Y(n6390) );
  INVX1 U3788 ( .A(fGx[3]), .Y(n6104) );
  NOR2X1 U3789 ( .A(n4048), .B(n5826), .Y(\U3/U122/Z_19 ) );
  INVX1 U3790 ( .A(fGx[20]), .Y(n4048) );
  NOR2X1 U3791 ( .A(n4046), .B(n5826), .Y(\U3/U122/Z_18 ) );
  INVX1 U3792 ( .A(fGx[19]), .Y(n4046) );
  NOR2X1 U3793 ( .A(n4044), .B(n5826), .Y(\U3/U122/Z_17 ) );
  INVX1 U3794 ( .A(fGx[18]), .Y(n4044) );
  NOR2X1 U3795 ( .A(n4042), .B(n5826), .Y(\U3/U122/Z_16 ) );
  INVX1 U3796 ( .A(fGx[17]), .Y(n4042) );
  NOR2X1 U3797 ( .A(n4040), .B(n5826), .Y(\U3/U122/Z_15 ) );
  INVX1 U3798 ( .A(fGx[16]), .Y(n4040) );
  NOR2X1 U3799 ( .A(n4038), .B(n5826), .Y(\U3/U122/Z_14 ) );
  INVX1 U3800 ( .A(fGx[15]), .Y(n4038) );
  NOR2X1 U3801 ( .A(n4036), .B(n5826), .Y(\U3/U122/Z_13 ) );
  INVX1 U3802 ( .A(fGx[14]), .Y(n4036) );
  NOR2X1 U3803 ( .A(n4034), .B(n5826), .Y(\U3/U122/Z_12 ) );
  INVX1 U3804 ( .A(fGx[13]), .Y(n4034) );
  NOR2X1 U3805 ( .A(n4032), .B(n5826), .Y(\U3/U122/Z_11 ) );
  INVX1 U3806 ( .A(fGx[12]), .Y(n4032) );
  NOR2X1 U3807 ( .A(n4030), .B(n5826), .Y(\U3/U122/Z_10 ) );
  INVX1 U3808 ( .A(fGx[11]), .Y(n4030) );
  OAI21X1 U3809 ( .A(n5826), .B(n6106), .C(n6391), .Y(\U3/U122/Z_1 ) );
  OAI21X1 U3810 ( .A(n6392), .B(n6393), .C(n7205), .Y(n6391) );
  NAND2X1 U3811 ( .A(n6394), .B(n6395), .Y(n6393) );
  NOR2X1 U3812 ( .A(n6396), .B(n6397), .Y(n6395) );
  OAI21X1 U3813 ( .A(n3830), .B(n6240), .C(n6398), .Y(n6397) );
  AOI22X1 U3814 ( .A(n6238), .B(\regX[1][1] ), .C(n6239), .D(\regX[11][1] ), 
        .Y(n6398) );
  INVX1 U3815 ( .A(\regX[7][1] ), .Y(n3830) );
  OAI21X1 U3816 ( .A(n3589), .B(n6258), .C(n6399), .Y(n6396) );
  AOI22X1 U3817 ( .A(n6242), .B(\regX[8][1] ), .C(n6243), .D(N1616), .Y(n6399)
         );
  INVX1 U3818 ( .A(\regX[23][1] ), .Y(n3589) );
  NOR2X1 U3819 ( .A(n6400), .B(n6401), .Y(n6394) );
  OAI21X1 U3820 ( .A(n3807), .B(n6236), .C(n6402), .Y(n6401) );
  AOI22X1 U3821 ( .A(n6352), .B(\regX[5][1] ), .C(n6353), .D(\regX[0][1] ), 
        .Y(n6402) );
  OAI21X1 U3822 ( .A(n3881), .B(n6320), .C(n6403), .Y(n6400) );
  AOI22X1 U3823 ( .A(n6228), .B(N1376), .C(n6233), .D(\regX[13][1] ), .Y(n6403) );
  INVX1 U3824 ( .A(N1434), .Y(n3881) );
  NAND3X1 U3825 ( .A(n6404), .B(n6405), .C(n6406), .Y(n6392) );
  NOR2X1 U3826 ( .A(n6407), .B(n6408), .Y(n6406) );
  OAI21X1 U3827 ( .A(n3655), .B(n6252), .C(n6409), .Y(n6408) );
  AOI22X1 U3828 ( .A(n6255), .B(\regX[15][1] ), .C(n6361), .D(N1678), .Y(n6409) );
  INVX1 U3829 ( .A(\regX[17][1] ), .Y(n3655) );
  OAI21X1 U3830 ( .A(n3634), .B(n6262), .C(n6410), .Y(n6407) );
  AOI22X1 U3831 ( .A(n6250), .B(\regX[16][1] ), .C(n6251), .D(N1736), .Y(n6410) );
  INVX1 U3832 ( .A(\regX[19][1] ), .Y(n3634) );
  NOR2X1 U3833 ( .A(n6411), .B(n6412), .Y(n6405) );
  OAI22X1 U3834 ( .A(n3602), .B(n6333), .C(n3624), .D(n6339), .Y(n6412) );
  INVX1 U3835 ( .A(\regX[20][1] ), .Y(n3624) );
  INVX1 U3836 ( .A(\regX[22][1] ), .Y(n3602) );
  OAI22X1 U3837 ( .A(n3563), .B(n6365), .C(n3843), .D(n6366), .Y(n6411) );
  INVX1 U3838 ( .A(\regX[24][1] ), .Y(n3563) );
  AOI21X1 U3839 ( .A(n6265), .B(\regX[18][1] ), .C(n6413), .Y(n6404) );
  OAI22X1 U3840 ( .A(n3613), .B(n6337), .C(n3893), .D(n6322), .Y(n6413) );
  INVX1 U3841 ( .A(\regX[3][1] ), .Y(n3893) );
  INVX1 U3842 ( .A(fGx[2]), .Y(n6106) );
  OAI21X1 U3843 ( .A(n5826), .B(n6108), .C(n6414), .Y(\U3/U122/Z_0 ) );
  OAI21X1 U3844 ( .A(n6415), .B(n6416), .C(n7205), .Y(n6414) );
  NAND2X1 U3845 ( .A(n6417), .B(n6418), .Y(n6416) );
  NOR2X1 U3846 ( .A(n6419), .B(n6420), .Y(n6418) );
  OAI21X1 U3847 ( .A(n3828), .B(n6240), .C(n6421), .Y(n6420) );
  AOI22X1 U3848 ( .A(n6238), .B(\regX[1][0] ), .C(n6239), .D(\regX[11][0] ), 
        .Y(n6421) );
  AND2X1 U3849 ( .A(n6422), .B(n6423), .Y(n6239) );
  AND2X1 U3850 ( .A(n6424), .B(n6425), .Y(n6238) );
  NAND2X1 U3851 ( .A(n6424), .B(n6426), .Y(n6240) );
  INVX1 U3852 ( .A(\regX[7][0] ), .Y(n3828) );
  OAI21X1 U3853 ( .A(n3587), .B(n6258), .C(n6427), .Y(n6419) );
  AOI22X1 U3854 ( .A(n6242), .B(\regX[8][0] ), .C(n6243), .D(N1615), .Y(n6427)
         );
  AND2X1 U3855 ( .A(n6422), .B(n6428), .Y(n6243) );
  INVX1 U3856 ( .A(n6429), .Y(n6242) );
  NAND3X1 U3857 ( .A(n6428), .B(n6425), .C(n6430), .Y(n6429) );
  NAND2X1 U3858 ( .A(n6431), .B(n6426), .Y(n6258) );
  INVX1 U3859 ( .A(\regX[23][0] ), .Y(n3587) );
  NOR2X1 U3860 ( .A(n6432), .B(n6433), .Y(n6417) );
  OAI21X1 U3861 ( .A(n3805), .B(n6236), .C(n6434), .Y(n6433) );
  AOI22X1 U3862 ( .A(n6352), .B(\regX[5][0] ), .C(n6353), .D(\regX[0][0] ), 
        .Y(n6434) );
  INVX1 U3863 ( .A(n6226), .Y(n6353) );
  NAND2X1 U3864 ( .A(n6435), .B(n6425), .Y(n6226) );
  INVX1 U3865 ( .A(n6230), .Y(n6352) );
  NAND2X1 U3866 ( .A(n6424), .B(n6436), .Y(n6230) );
  NAND2X1 U3867 ( .A(n6425), .B(n6423), .Y(n6236) );
  OAI21X1 U3868 ( .A(n3879), .B(n6320), .C(n6437), .Y(n6432) );
  AOI22X1 U3869 ( .A(n6228), .B(N1375), .C(n6233), .D(\regX[13][0] ), .Y(n6437) );
  AND2X1 U3870 ( .A(n6436), .B(n6423), .Y(n6233) );
  AND2X1 U3871 ( .A(n6435), .B(n6422), .Y(n6228) );
  NAND2X1 U3872 ( .A(n6435), .B(n6436), .Y(n6320) );
  INVX1 U3873 ( .A(N1433), .Y(n3879) );
  NAND3X1 U3874 ( .A(n6438), .B(n6439), .C(n6440), .Y(n6415) );
  NOR2X1 U3875 ( .A(n6441), .B(n6442), .Y(n6440) );
  OAI21X1 U3876 ( .A(n3653), .B(n6252), .C(n6443), .Y(n6442) );
  AOI22X1 U3877 ( .A(n6255), .B(\regX[15][0] ), .C(n6361), .D(N1677), .Y(n6443) );
  INVX1 U3878 ( .A(n6248), .Y(n6361) );
  NAND2X1 U3879 ( .A(n6436), .B(n6428), .Y(n6248) );
  AND2X1 U3880 ( .A(n6423), .B(n6426), .Y(n6255) );
  NOR2X1 U3881 ( .A(n6444), .B(n6445), .Y(n6423) );
  NAND2X1 U3882 ( .A(n6425), .B(n6431), .Y(n6252) );
  INVX1 U3883 ( .A(\regX[17][0] ), .Y(n3653) );
  OAI21X1 U3884 ( .A(n3632), .B(n6262), .C(n6446), .Y(n6441) );
  AOI22X1 U3885 ( .A(n6250), .B(\regX[16][0] ), .C(n6251), .D(N1735), .Y(n6446) );
  AND2X1 U3886 ( .A(n6428), .B(n6426), .Y(n6251) );
  NOR2X1 U3887 ( .A(n6444), .B(n6447), .Y(n6428) );
  INVX1 U3888 ( .A(n6448), .Y(n6250) );
  NAND3X1 U3889 ( .A(n6449), .B(n6444), .C(n6425), .Y(n6448) );
  NOR2X1 U3890 ( .A(n6450), .B(n6451), .Y(n6425) );
  NAND2X1 U3891 ( .A(n6422), .B(n6431), .Y(n6262) );
  INVX1 U3892 ( .A(\regX[19][0] ), .Y(n3632) );
  NOR2X1 U3893 ( .A(n6452), .B(n6453), .Y(n6439) );
  OAI22X1 U3894 ( .A(n3600), .B(n6333), .C(n3622), .D(n6339), .Y(n6453) );
  NAND2X1 U3895 ( .A(n6436), .B(n6449), .Y(n6339) );
  NAND2X1 U3896 ( .A(n6426), .B(n6449), .Y(n6333) );
  OAI22X1 U3897 ( .A(n3560), .B(n6365), .C(n3841), .D(n6366), .Y(n6452) );
  NAND2X1 U3898 ( .A(n6435), .B(n6426), .Y(n6366) );
  NOR2X1 U3899 ( .A(n6454), .B(n6455), .Y(n6426) );
  INVX1 U3900 ( .A(n6456), .Y(n6435) );
  NAND3X1 U3901 ( .A(n6445), .B(n6444), .C(n6430), .Y(n6456) );
  INVX1 U3902 ( .A(n6260), .Y(n6365) );
  NOR2X1 U3903 ( .A(n6444), .B(n6430), .Y(n6260) );
  AOI21X1 U3904 ( .A(n6265), .B(\regX[18][0] ), .C(n6457), .Y(n6438) );
  OAI22X1 U3905 ( .A(n3611), .B(n6337), .C(n3891), .D(n6322), .Y(n6457) );
  NAND2X1 U3906 ( .A(n6424), .B(n6422), .Y(n6322) );
  INVX1 U3907 ( .A(n6458), .Y(n6424) );
  NAND3X1 U3908 ( .A(n6444), .B(n6447), .C(n6430), .Y(n6458) );
  NAND2X1 U3909 ( .A(n6436), .B(n6431), .Y(n6337) );
  NOR2X1 U3910 ( .A(n6445), .B(n6430), .Y(n6431) );
  NOR2X1 U3911 ( .A(n6455), .B(n6451), .Y(n6436) );
  INVX1 U3912 ( .A(n6450), .Y(n6455) );
  AND2X1 U3913 ( .A(n6422), .B(n6449), .Y(n6265) );
  NOR2X1 U3914 ( .A(n6447), .B(n6430), .Y(n6449) );
  XNOR2X1 U3915 ( .A(n6459), .B(n6460), .Y(n6430) );
  XOR2X1 U3916 ( .A(n6461), .B(n6066), .Y(n6459) );
  XNOR2X1 U3917 ( .A(n6462), .B(n6463), .Y(n6066) );
  AOI21X1 U3918 ( .A(n7246), .B(N3093), .C(n6464), .Y(n6463) );
  OAI21X1 U3919 ( .A(n6465), .B(n6466), .C(n6467), .Y(n6462) );
  OAI21X1 U3920 ( .A(n6468), .B(n6469), .C(n6470), .Y(n6467) );
  OAI21X1 U3921 ( .A(n6471), .B(n6472), .C(n6473), .Y(n6461) );
  OAI21X1 U3922 ( .A(n6474), .B(n6475), .C(n6476), .Y(n6473) );
  INVX1 U3923 ( .A(n6472), .Y(n6474) );
  NOR2X1 U3924 ( .A(n6454), .B(n6450), .Y(n6422) );
  XOR2X1 U3925 ( .A(n6477), .B(n6476), .Y(n6450) );
  XOR2X1 U3926 ( .A(n6075), .B(n6478), .Y(n6477) );
  INVX1 U3927 ( .A(fGx[1]), .Y(n6108) );
  AND2X1 U3928 ( .A(fGy[7]), .B(n7240), .Y(\U3/U121/Z_7 ) );
  AND2X1 U3929 ( .A(fGy[6]), .B(n7240), .Y(\U3/U121/Z_6 ) );
  AND2X1 U3930 ( .A(fGy[5]), .B(n7240), .Y(\U3/U121/Z_5 ) );
  AND2X1 U3931 ( .A(fGy[4]), .B(n7240), .Y(\U3/U121/Z_4 ) );
  OAI21X1 U3932 ( .A(n5826), .B(n6479), .C(n6480), .Y(\U3/U121/Z_3 ) );
  OAI21X1 U3933 ( .A(n5826), .B(n6481), .C(n6480), .Y(\U3/U121/Z_2 ) );
  INVX1 U3934 ( .A(fGy[2]), .Y(n6481) );
  OAI21X1 U3935 ( .A(n5826), .B(n6482), .C(n6480), .Y(\U3/U121/Z_1 ) );
  OAI21X1 U3936 ( .A(n5826), .B(n6483), .C(n6480), .Y(\U3/U121/Z_0 ) );
  INVX1 U3937 ( .A(fGy[0]), .Y(n6483) );
  NAND2X1 U3938 ( .A(n4080), .B(n3467), .Y(n5826) );
  NOR2X1 U3939 ( .A(n3477), .B(n6200), .Y(\U3/U119/Z_9 ) );
  INVX1 U3940 ( .A(N2755), .Y(n6200) );
  NOR2X1 U3941 ( .A(n3477), .B(n6175), .Y(\U3/U119/Z_8 ) );
  INVX1 U3942 ( .A(N2754), .Y(n6175) );
  NAND3X1 U3943 ( .A(n6484), .B(n6485), .C(n6486), .Y(\U3/U119/Z_7 ) );
  NOR2X1 U3944 ( .A(n6487), .B(n6488), .Y(n6486) );
  OR2X1 U3945 ( .A(n6489), .B(n6490), .Y(n6488) );
  OAI21X1 U3946 ( .A(n3661), .B(n6491), .C(n6492), .Y(n6490) );
  AOI22X1 U3947 ( .A(n6493), .B(\regX[16][7] ), .C(n6494), .D(\regX[24][7] ), 
        .Y(n6492) );
  INVX1 U3948 ( .A(\regX[17][7] ), .Y(n3661) );
  OAI21X1 U3949 ( .A(n3887), .B(n6495), .C(n6496), .Y(n6489) );
  AOI22X1 U3950 ( .A(n6497), .B(\regX[15][7] ), .C(n6498), .D(N1742), .Y(n6496) );
  INVX1 U3951 ( .A(N1440), .Y(n3887) );
  NAND3X1 U3952 ( .A(n6499), .B(n6500), .C(n6501), .Y(n6487) );
  AOI21X1 U3953 ( .A(n6502), .B(\regX[21][7] ), .C(n6503), .Y(n6501) );
  OAI22X1 U3954 ( .A(n3595), .B(n6504), .C(n3651), .D(n6505), .Y(n6503) );
  INVX1 U3955 ( .A(\regX[23][7] ), .Y(n3595) );
  AOI22X1 U3956 ( .A(n6506), .B(N1684), .C(n6507), .D(\regX[19][7] ), .Y(n6500) );
  AOI22X1 U3957 ( .A(n6508), .B(\regX[13][7] ), .C(n6509), .D(\regX[20][7] ), 
        .Y(n6499) );
  NOR2X1 U3958 ( .A(n6510), .B(n6511), .Y(n6485) );
  OAI21X1 U3959 ( .A(n3932), .B(n6512), .C(n6513), .Y(n6511) );
  AOI22X1 U3960 ( .A(n6514), .B(\regX[22][7] ), .C(n6515), .D(\regX[1][7] ), 
        .Y(n6513) );
  INVX1 U3961 ( .A(\regX[0][7] ), .Y(n3932) );
  OR2X1 U3962 ( .A(n6516), .B(n6517), .Y(n6510) );
  OAI22X1 U3963 ( .A(n3825), .B(n6518), .C(n3813), .D(n6519), .Y(n6517) );
  OAI21X1 U3964 ( .A(n3836), .B(n6520), .C(n3525), .Y(n6516) );
  NAND2X1 U3965 ( .A(N2753), .B(n3467), .Y(n3525) );
  INVX1 U3966 ( .A(\regX[7][7] ), .Y(n3836) );
  NOR2X1 U3967 ( .A(n6521), .B(n6522), .Y(n6484) );
  OAI21X1 U3968 ( .A(n3899), .B(n6523), .C(n6524), .Y(n6522) );
  AOI22X1 U3969 ( .A(n6525), .B(N1382), .C(\regX[6][7] ), .D(n6526), .Y(n6524)
         );
  OAI21X1 U3970 ( .A(n3794), .B(n6527), .C(n6528), .Y(n6521) );
  AOI22X1 U3971 ( .A(n6529), .B(\regX[5][7] ), .C(n6530), .D(N1622), .Y(n6528)
         );
  INVX1 U3972 ( .A(\regX[11][7] ), .Y(n3794) );
  NAND3X1 U3973 ( .A(n6531), .B(n6532), .C(n6533), .Y(\U3/U119/Z_6 ) );
  NOR2X1 U3974 ( .A(n6534), .B(n6535), .Y(n6533) );
  OR2X1 U3975 ( .A(n6536), .B(n6537), .Y(n6535) );
  OAI21X1 U3976 ( .A(n3660), .B(n6491), .C(n6538), .Y(n6537) );
  AOI22X1 U3977 ( .A(n6493), .B(\regX[16][6] ), .C(n6494), .D(\regX[24][6] ), 
        .Y(n6538) );
  INVX1 U3978 ( .A(\regX[17][6] ), .Y(n3660) );
  OAI21X1 U3979 ( .A(n3886), .B(n6495), .C(n6539), .Y(n6536) );
  AOI22X1 U3980 ( .A(n6497), .B(\regX[15][6] ), .C(n6498), .D(N1741), .Y(n6539) );
  INVX1 U3981 ( .A(N1439), .Y(n3886) );
  NAND3X1 U3982 ( .A(n6540), .B(n6541), .C(n6542), .Y(n6534) );
  AOI21X1 U3983 ( .A(n6502), .B(\regX[21][6] ), .C(n6543), .Y(n6542) );
  OAI22X1 U3984 ( .A(n3594), .B(n6504), .C(n3650), .D(n6505), .Y(n6543) );
  INVX1 U3985 ( .A(\regX[23][6] ), .Y(n3594) );
  AOI22X1 U3986 ( .A(n6506), .B(N1683), .C(n6507), .D(\regX[19][6] ), .Y(n6541) );
  AOI22X1 U3987 ( .A(n6508), .B(\regX[13][6] ), .C(n6509), .D(\regX[20][6] ), 
        .Y(n6540) );
  NOR2X1 U3988 ( .A(n6544), .B(n6545), .Y(n6532) );
  OAI21X1 U3989 ( .A(n3931), .B(n6512), .C(n6546), .Y(n6545) );
  AOI22X1 U3990 ( .A(n6514), .B(\regX[22][6] ), .C(n6515), .D(\regX[1][6] ), 
        .Y(n6546) );
  INVX1 U3991 ( .A(\regX[0][6] ), .Y(n3931) );
  OR2X1 U3992 ( .A(n6547), .B(n6548), .Y(n6544) );
  OAI22X1 U3993 ( .A(n3824), .B(n6518), .C(n3812), .D(n6519), .Y(n6548) );
  OAI21X1 U3994 ( .A(n3835), .B(n6520), .C(n3526), .Y(n6547) );
  NAND2X1 U3995 ( .A(N2752), .B(n3467), .Y(n3526) );
  INVX1 U3996 ( .A(\regX[7][6] ), .Y(n3835) );
  NOR2X1 U3997 ( .A(n6549), .B(n6550), .Y(n6531) );
  OAI21X1 U3998 ( .A(n3898), .B(n6523), .C(n6551), .Y(n6550) );
  AOI22X1 U3999 ( .A(n6525), .B(N1381), .C(\regX[6][6] ), .D(n6526), .Y(n6551)
         );
  OAI21X1 U4000 ( .A(n3793), .B(n6527), .C(n6552), .Y(n6549) );
  AOI22X1 U4001 ( .A(n6529), .B(\regX[5][6] ), .C(n6530), .D(N1621), .Y(n6552)
         );
  INVX1 U4002 ( .A(\regX[11][6] ), .Y(n3793) );
  NAND3X1 U4003 ( .A(n6553), .B(n6554), .C(n6555), .Y(\U3/U119/Z_5 ) );
  NOR2X1 U4004 ( .A(n6556), .B(n6557), .Y(n6555) );
  OR2X1 U4005 ( .A(n6558), .B(n6559), .Y(n6557) );
  OAI21X1 U4006 ( .A(n3659), .B(n6491), .C(n6560), .Y(n6559) );
  AOI22X1 U4007 ( .A(n6493), .B(\regX[16][5] ), .C(n6494), .D(\regX[24][5] ), 
        .Y(n6560) );
  INVX1 U4008 ( .A(\regX[17][5] ), .Y(n3659) );
  OAI21X1 U4009 ( .A(n3885), .B(n6495), .C(n6561), .Y(n6558) );
  AOI22X1 U4010 ( .A(n6497), .B(\regX[15][5] ), .C(n6498), .D(N1740), .Y(n6561) );
  INVX1 U4011 ( .A(N1438), .Y(n3885) );
  NAND3X1 U4012 ( .A(n6562), .B(n6563), .C(n6564), .Y(n6556) );
  AOI21X1 U4013 ( .A(n6502), .B(\regX[21][5] ), .C(n6565), .Y(n6564) );
  OAI22X1 U4014 ( .A(n3593), .B(n6504), .C(n3649), .D(n6505), .Y(n6565) );
  INVX1 U4015 ( .A(\regX[23][5] ), .Y(n3593) );
  AOI22X1 U4016 ( .A(n6506), .B(N1682), .C(n6507), .D(\regX[19][5] ), .Y(n6563) );
  AOI22X1 U4017 ( .A(n6508), .B(\regX[13][5] ), .C(n6509), .D(\regX[20][5] ), 
        .Y(n6562) );
  NOR2X1 U4018 ( .A(n6566), .B(n6567), .Y(n6554) );
  OAI21X1 U4019 ( .A(n3930), .B(n6512), .C(n6568), .Y(n6567) );
  AOI22X1 U4020 ( .A(n6514), .B(\regX[22][5] ), .C(n6515), .D(\regX[1][5] ), 
        .Y(n6568) );
  INVX1 U4021 ( .A(\regX[0][5] ), .Y(n3930) );
  OR2X1 U4022 ( .A(n6569), .B(n6570), .Y(n6566) );
  OAI22X1 U4023 ( .A(n3823), .B(n6518), .C(n3811), .D(n6519), .Y(n6570) );
  OAI21X1 U4024 ( .A(n3834), .B(n6520), .C(n3527), .Y(n6569) );
  NAND2X1 U4025 ( .A(N2751), .B(n3467), .Y(n3527) );
  INVX1 U4026 ( .A(\regX[7][5] ), .Y(n3834) );
  NOR2X1 U4027 ( .A(n6571), .B(n6572), .Y(n6553) );
  OAI21X1 U4028 ( .A(n3897), .B(n6523), .C(n6573), .Y(n6572) );
  AOI22X1 U4029 ( .A(n6525), .B(N1380), .C(\regX[6][5] ), .D(n6526), .Y(n6573)
         );
  OAI21X1 U4030 ( .A(n3792), .B(n6527), .C(n6574), .Y(n6571) );
  AOI22X1 U4031 ( .A(n6529), .B(\regX[5][5] ), .C(n6530), .D(N1620), .Y(n6574)
         );
  INVX1 U4032 ( .A(\regX[11][5] ), .Y(n3792) );
  NAND3X1 U4033 ( .A(n6575), .B(n6576), .C(n6577), .Y(\U3/U119/Z_4 ) );
  NOR2X1 U4034 ( .A(n6578), .B(n6579), .Y(n6577) );
  OR2X1 U4035 ( .A(n6580), .B(n6581), .Y(n6579) );
  OAI21X1 U4036 ( .A(n3658), .B(n6491), .C(n6582), .Y(n6581) );
  AOI22X1 U4037 ( .A(n6493), .B(\regX[16][4] ), .C(n6494), .D(\regX[24][4] ), 
        .Y(n6582) );
  INVX1 U4038 ( .A(n6583), .Y(n6493) );
  INVX1 U4039 ( .A(\regX[17][4] ), .Y(n3658) );
  OAI21X1 U4040 ( .A(n3884), .B(n6495), .C(n6584), .Y(n6580) );
  AOI22X1 U4041 ( .A(n6497), .B(\regX[15][4] ), .C(n6498), .D(N1739), .Y(n6584) );
  INVX1 U4042 ( .A(N1437), .Y(n3884) );
  NAND3X1 U4043 ( .A(n6585), .B(n6586), .C(n6587), .Y(n6578) );
  AOI21X1 U4044 ( .A(n6502), .B(\regX[21][4] ), .C(n6588), .Y(n6587) );
  OAI22X1 U4045 ( .A(n3592), .B(n6504), .C(n3648), .D(n6505), .Y(n6588) );
  INVX1 U4046 ( .A(n6589), .Y(n6504) );
  INVX1 U4047 ( .A(\regX[23][4] ), .Y(n3592) );
  AOI22X1 U4048 ( .A(n6506), .B(N1681), .C(n6507), .D(\regX[19][4] ), .Y(n6586) );
  INVX1 U4049 ( .A(n6590), .Y(n6506) );
  AOI22X1 U4050 ( .A(n6508), .B(\regX[13][4] ), .C(n6509), .D(\regX[20][4] ), 
        .Y(n6585) );
  NOR2X1 U4051 ( .A(n6591), .B(n6592), .Y(n6576) );
  OAI21X1 U4052 ( .A(n3929), .B(n6512), .C(n6593), .Y(n6592) );
  AOI22X1 U4053 ( .A(n6514), .B(\regX[22][4] ), .C(n6515), .D(\regX[1][4] ), 
        .Y(n6593) );
  INVX1 U4054 ( .A(n6594), .Y(n6515) );
  INVX1 U4055 ( .A(\regX[0][4] ), .Y(n3929) );
  OR2X1 U4056 ( .A(n6595), .B(n6596), .Y(n6591) );
  OAI22X1 U4057 ( .A(n3822), .B(n6518), .C(n3810), .D(n6519), .Y(n6596) );
  OAI21X1 U4058 ( .A(n3833), .B(n6520), .C(n3528), .Y(n6595) );
  NAND2X1 U4059 ( .A(N2750), .B(n3467), .Y(n3528) );
  INVX1 U4060 ( .A(n6597), .Y(n6520) );
  INVX1 U4061 ( .A(\regX[7][4] ), .Y(n3833) );
  NOR2X1 U4062 ( .A(n6598), .B(n6599), .Y(n6575) );
  OAI21X1 U4063 ( .A(n3896), .B(n6523), .C(n6600), .Y(n6599) );
  AOI22X1 U4064 ( .A(n6525), .B(N1379), .C(\regX[6][4] ), .D(n6526), .Y(n6600)
         );
  INVX1 U4065 ( .A(n6601), .Y(n6525) );
  OAI21X1 U4066 ( .A(n3791), .B(n6527), .C(n6602), .Y(n6598) );
  AOI22X1 U4067 ( .A(n6529), .B(\regX[5][4] ), .C(n6530), .D(N1619), .Y(n6602)
         );
  INVX1 U4068 ( .A(\regX[11][4] ), .Y(n3791) );
  NOR2X1 U4069 ( .A(n3477), .B(n6177), .Y(\U3/U119/Z_31 ) );
  INVX1 U4070 ( .A(N2776), .Y(n6177) );
  NAND3X1 U4071 ( .A(n6603), .B(n6604), .C(n6605), .Y(\U3/U119/Z_3 ) );
  NOR2X1 U4072 ( .A(n6606), .B(n6607), .Y(n6605) );
  OR2X1 U4073 ( .A(n6608), .B(n6609), .Y(n6607) );
  OAI21X1 U4074 ( .A(n3780), .B(n6590), .C(n6610), .Y(n6609) );
  AOI22X1 U4075 ( .A(\regX[6][3] ), .B(n6526), .C(n6611), .D(\regX[3][3] ), 
        .Y(n6610) );
  OAI21X1 U4076 ( .A(n3907), .B(n6601), .C(n6612), .Y(n6608) );
  AOI22X1 U4077 ( .A(n6530), .B(N1618), .C(n6613), .D(\regX[11][3] ), .Y(n6612) );
  NAND3X1 U4078 ( .A(n6614), .B(n6615), .C(n6616), .Y(n6606) );
  AOI21X1 U4079 ( .A(n6529), .B(\regX[5][3] ), .C(n6617), .Y(n6616) );
  OAI22X1 U4080 ( .A(n3928), .B(n6512), .C(n3918), .D(n6594), .Y(n6617) );
  INVX1 U4081 ( .A(\regX[0][3] ), .Y(n3928) );
  AOI22X1 U4082 ( .A(n6597), .B(\regX[7][3] ), .C(n6618), .D(\regX[9][3] ), 
        .Y(n6615) );
  AOI22X1 U4083 ( .A(n6619), .B(\regX[8][3] ), .C(n6514), .D(\regX[22][3] ), 
        .Y(n6614) );
  NOR2X1 U4084 ( .A(n6620), .B(n6621), .Y(n6604) );
  OAI21X1 U4085 ( .A(n3749), .B(n6622), .C(n6623), .Y(n6621) );
  AOI22X1 U4086 ( .A(n6589), .B(\regX[23][3] ), .C(n6502), .D(\regX[21][3] ), 
        .Y(n6623) );
  NAND2X1 U4087 ( .A(n6624), .B(n6625), .Y(n6620) );
  AOI22X1 U4088 ( .A(n6507), .B(\regX[19][3] ), .C(n6508), .D(\regX[13][3] ), 
        .Y(n6625) );
  AOI22X1 U4089 ( .A(n6509), .B(\regX[20][3] ), .C(n6626), .D(\regX[18][3] ), 
        .Y(n6624) );
  NOR2X1 U4090 ( .A(n6627), .B(n6628), .Y(n6603) );
  OAI21X1 U4091 ( .A(n3477), .B(n6176), .C(n6629), .Y(n6628) );
  AOI22X1 U4092 ( .A(n6494), .B(\regX[24][3] ), .C(n6630), .D(\regX[17][3] ), 
        .Y(n6629) );
  OAI21X1 U4093 ( .A(n3670), .B(n6583), .C(n6631), .Y(n6627) );
  AOI22X1 U4094 ( .A(n6498), .B(N1738), .C(n6632), .D(N1436), .Y(n6631) );
  INVX1 U4095 ( .A(\regX[16][3] ), .Y(n3670) );
  NOR2X1 U4096 ( .A(n3477), .B(n6178), .Y(\U3/U119/Z_29 ) );
  INVX1 U4097 ( .A(N2775), .Y(n6178) );
  NOR2X1 U4098 ( .A(n3477), .B(n6180), .Y(\U3/U119/Z_28 ) );
  INVX1 U4099 ( .A(N2774), .Y(n6180) );
  NOR2X1 U4100 ( .A(n3477), .B(n6181), .Y(\U3/U119/Z_27 ) );
  INVX1 U4101 ( .A(N2773), .Y(n6181) );
  NOR2X1 U4102 ( .A(n3477), .B(n6182), .Y(\U3/U119/Z_26 ) );
  INVX1 U4103 ( .A(N2772), .Y(n6182) );
  NOR2X1 U4104 ( .A(n3477), .B(n6183), .Y(\U3/U119/Z_25 ) );
  INVX1 U4105 ( .A(N2771), .Y(n6183) );
  NOR2X1 U4106 ( .A(n3477), .B(n6184), .Y(\U3/U119/Z_24 ) );
  INVX1 U4107 ( .A(N2770), .Y(n6184) );
  NOR2X1 U4108 ( .A(n3477), .B(n6185), .Y(\U3/U119/Z_23 ) );
  INVX1 U4109 ( .A(N2769), .Y(n6185) );
  NOR2X1 U4110 ( .A(n3477), .B(n6186), .Y(\U3/U119/Z_22 ) );
  INVX1 U4111 ( .A(N2768), .Y(n6186) );
  NOR2X1 U4112 ( .A(n3477), .B(n6187), .Y(\U3/U119/Z_21 ) );
  INVX1 U4113 ( .A(N2767), .Y(n6187) );
  NOR2X1 U4114 ( .A(n3477), .B(n6188), .Y(\U3/U119/Z_20 ) );
  INVX1 U4115 ( .A(N2766), .Y(n6188) );
  NAND3X1 U4116 ( .A(n6633), .B(n6634), .C(n6635), .Y(\U3/U119/Z_2 ) );
  NOR2X1 U4117 ( .A(n6636), .B(n6637), .Y(n6635) );
  OR2X1 U4118 ( .A(n6638), .B(n6639), .Y(n6637) );
  OAI21X1 U4119 ( .A(n3779), .B(n6590), .C(n6640), .Y(n6639) );
  AOI22X1 U4120 ( .A(\regX[6][2] ), .B(n6526), .C(n6611), .D(\regX[3][2] ), 
        .Y(n6640) );
  OAI21X1 U4121 ( .A(n3906), .B(n6601), .C(n6641), .Y(n6638) );
  AOI22X1 U4122 ( .A(n6530), .B(N1617), .C(n6613), .D(\regX[11][2] ), .Y(n6641) );
  NAND3X1 U4123 ( .A(n6642), .B(n6643), .C(n6644), .Y(n6636) );
  AOI21X1 U4124 ( .A(n6529), .B(\regX[5][2] ), .C(n6645), .Y(n6644) );
  OAI22X1 U4125 ( .A(n3926), .B(n6512), .C(n3917), .D(n6594), .Y(n6645) );
  INVX1 U4126 ( .A(\regX[0][2] ), .Y(n3926) );
  AOI22X1 U4127 ( .A(n6597), .B(\regX[7][2] ), .C(n6618), .D(\regX[9][2] ), 
        .Y(n6643) );
  AOI22X1 U4128 ( .A(n6619), .B(\regX[8][2] ), .C(n6514), .D(\regX[22][2] ), 
        .Y(n6642) );
  NOR2X1 U4129 ( .A(n6646), .B(n6647), .Y(n6634) );
  OAI21X1 U4130 ( .A(n3740), .B(n6622), .C(n6648), .Y(n6647) );
  AOI22X1 U4131 ( .A(n6589), .B(\regX[23][2] ), .C(n6502), .D(\regX[21][2] ), 
        .Y(n6648) );
  NAND2X1 U4132 ( .A(n6649), .B(n6650), .Y(n6646) );
  AOI22X1 U4133 ( .A(n6507), .B(\regX[19][2] ), .C(n6508), .D(\regX[13][2] ), 
        .Y(n6650) );
  AOI22X1 U4134 ( .A(n6509), .B(\regX[20][2] ), .C(n6626), .D(\regX[18][2] ), 
        .Y(n6649) );
  NOR2X1 U4135 ( .A(n6651), .B(n6652), .Y(n6633) );
  OAI21X1 U4136 ( .A(n3477), .B(n6179), .C(n6653), .Y(n6652) );
  AOI22X1 U4137 ( .A(n6494), .B(\regX[24][2] ), .C(n6630), .D(\regX[17][2] ), 
        .Y(n6653) );
  OAI21X1 U4138 ( .A(n3669), .B(n6583), .C(n6654), .Y(n6651) );
  AOI22X1 U4139 ( .A(n6498), .B(N1737), .C(n6632), .D(N1435), .Y(n6654) );
  INVX1 U4140 ( .A(\regX[16][2] ), .Y(n3669) );
  NOR2X1 U4141 ( .A(n3477), .B(n6189), .Y(\U3/U119/Z_19 ) );
  INVX1 U4142 ( .A(N2765), .Y(n6189) );
  NOR2X1 U4143 ( .A(n3477), .B(n6191), .Y(\U3/U119/Z_18 ) );
  INVX1 U4144 ( .A(N2764), .Y(n6191) );
  NOR2X1 U4145 ( .A(n3477), .B(n6192), .Y(\U3/U119/Z_17 ) );
  INVX1 U4146 ( .A(N2763), .Y(n6192) );
  NOR2X1 U4147 ( .A(n3477), .B(n6193), .Y(\U3/U119/Z_16 ) );
  INVX1 U4148 ( .A(N2762), .Y(n6193) );
  NOR2X1 U4149 ( .A(n3477), .B(n6194), .Y(\U3/U119/Z_15 ) );
  INVX1 U4150 ( .A(N2761), .Y(n6194) );
  NOR2X1 U4151 ( .A(n3477), .B(n6195), .Y(\U3/U119/Z_14 ) );
  INVX1 U4152 ( .A(N2760), .Y(n6195) );
  NOR2X1 U4153 ( .A(n3477), .B(n6196), .Y(\U3/U119/Z_13 ) );
  INVX1 U4154 ( .A(N2759), .Y(n6196) );
  NOR2X1 U4155 ( .A(n3477), .B(n6197), .Y(\U3/U119/Z_12 ) );
  INVX1 U4156 ( .A(N2758), .Y(n6197) );
  NOR2X1 U4157 ( .A(n3477), .B(n6198), .Y(\U3/U119/Z_11 ) );
  INVX1 U4158 ( .A(N2757), .Y(n6198) );
  NOR2X1 U4159 ( .A(n3477), .B(n6199), .Y(\U3/U119/Z_10 ) );
  INVX1 U4160 ( .A(N2756), .Y(n6199) );
  NAND3X1 U4161 ( .A(n6655), .B(n6656), .C(n6657), .Y(\U3/U119/Z_1 ) );
  NOR2X1 U4162 ( .A(n6658), .B(n6659), .Y(n6657) );
  OR2X1 U4163 ( .A(n6660), .B(n6661), .Y(n6659) );
  OAI21X1 U4164 ( .A(n3778), .B(n6590), .C(n6662), .Y(n6661) );
  AOI22X1 U4165 ( .A(\regX[6][1] ), .B(n6526), .C(n6611), .D(\regX[3][1] ), 
        .Y(n6662) );
  OAI21X1 U4166 ( .A(n3905), .B(n6601), .C(n6663), .Y(n6660) );
  AOI22X1 U4167 ( .A(n6530), .B(N1616), .C(n6613), .D(\regX[11][1] ), .Y(n6663) );
  NAND3X1 U4168 ( .A(n6664), .B(n6665), .C(n6666), .Y(n6658) );
  AOI21X1 U4169 ( .A(n6529), .B(\regX[5][1] ), .C(n6667), .Y(n6666) );
  OAI22X1 U4170 ( .A(n3934), .B(n6512), .C(n3916), .D(n6594), .Y(n6667) );
  INVX1 U4171 ( .A(\regX[0][1] ), .Y(n3934) );
  AOI22X1 U4172 ( .A(n6597), .B(\regX[7][1] ), .C(n6618), .D(\regX[9][1] ), 
        .Y(n6665) );
  AOI22X1 U4173 ( .A(n6619), .B(\regX[8][1] ), .C(n6514), .D(\regX[22][1] ), 
        .Y(n6664) );
  NOR2X1 U4174 ( .A(n6668), .B(n6669), .Y(n6656) );
  OAI21X1 U4175 ( .A(n3681), .B(n6622), .C(n6670), .Y(n6669) );
  AOI22X1 U4176 ( .A(n6589), .B(\regX[23][1] ), .C(n6502), .D(\regX[21][1] ), 
        .Y(n6670) );
  NAND2X1 U4177 ( .A(n6671), .B(n6672), .Y(n6668) );
  AOI22X1 U4178 ( .A(n6507), .B(\regX[19][1] ), .C(n6508), .D(\regX[13][1] ), 
        .Y(n6672) );
  AOI22X1 U4179 ( .A(n6509), .B(\regX[20][1] ), .C(n6626), .D(\regX[18][1] ), 
        .Y(n6671) );
  NOR2X1 U4180 ( .A(n6673), .B(n6674), .Y(n6655) );
  OAI21X1 U4181 ( .A(n3477), .B(n6190), .C(n6675), .Y(n6674) );
  AOI22X1 U4182 ( .A(n6494), .B(\regX[24][1] ), .C(n6630), .D(\regX[17][1] ), 
        .Y(n6675) );
  OAI21X1 U4183 ( .A(n3668), .B(n6583), .C(n6676), .Y(n6673) );
  AOI22X1 U4184 ( .A(n6498), .B(N1736), .C(n6632), .D(N1434), .Y(n6676) );
  INVX1 U4185 ( .A(\regX[16][1] ), .Y(n3668) );
  NAND3X1 U4186 ( .A(n6677), .B(n6678), .C(n6679), .Y(\U3/U119/Z_0 ) );
  NOR2X1 U4187 ( .A(n6680), .B(n6681), .Y(n6679) );
  OR2X1 U4188 ( .A(n6682), .B(n6683), .Y(n6681) );
  OAI21X1 U4189 ( .A(n3776), .B(n6590), .C(n6684), .Y(n6683) );
  AOI22X1 U4190 ( .A(\regX[6][0] ), .B(n6526), .C(n6611), .D(\regX[3][0] ), 
        .Y(n6684) );
  INVX1 U4191 ( .A(n6523), .Y(n6611) );
  NAND2X1 U4192 ( .A(n6685), .B(n6686), .Y(n6523) );
  OAI21X1 U4193 ( .A(n6687), .B(n6688), .C(n5827), .Y(n6526) );
  NAND2X1 U4194 ( .A(n6689), .B(n6690), .Y(n6590) );
  INVX1 U4195 ( .A(N1677), .Y(n3776) );
  OAI21X1 U4196 ( .A(n3903), .B(n6601), .C(n6691), .Y(n6682) );
  AOI22X1 U4197 ( .A(n6530), .B(N1615), .C(n6613), .D(\regX[11][0] ), .Y(n6691) );
  INVX1 U4198 ( .A(n6527), .Y(n6613) );
  NAND2X1 U4199 ( .A(n6685), .B(n6692), .Y(n6527) );
  AND2X1 U4200 ( .A(n6685), .B(n6690), .Y(n6530) );
  NAND2X1 U4201 ( .A(n6685), .B(n6693), .Y(n6601) );
  NAND3X1 U4202 ( .A(n6694), .B(n6695), .C(n6696), .Y(n6680) );
  AOI21X1 U4203 ( .A(n6529), .B(\regX[5][0] ), .C(n6697), .Y(n6696) );
  OAI22X1 U4204 ( .A(n3933), .B(n6512), .C(n3914), .D(n6594), .Y(n6697) );
  NAND2X1 U4205 ( .A(n6698), .B(n6686), .Y(n6594) );
  NAND2X1 U4206 ( .A(n6693), .B(n6698), .Y(n6512) );
  INVX1 U4207 ( .A(\regX[0][0] ), .Y(n3933) );
  AND2X1 U4208 ( .A(n6689), .B(n6686), .Y(n6529) );
  INVX1 U4209 ( .A(n6699), .Y(n6686) );
  AOI22X1 U4210 ( .A(n6597), .B(\regX[7][0] ), .C(n6618), .D(\regX[9][0] ), 
        .Y(n6695) );
  INVX1 U4211 ( .A(n6519), .Y(n6618) );
  NAND2X1 U4212 ( .A(n6698), .B(n6692), .Y(n6519) );
  NOR2X1 U4213 ( .A(n6687), .B(n6699), .Y(n6597) );
  NAND3X1 U4214 ( .A(n6700), .B(n6701), .C(n6702), .Y(n6699) );
  NOR2X1 U4215 ( .A(n6480), .B(n6703), .Y(n6702) );
  AOI22X1 U4216 ( .A(n6619), .B(\regX[8][0] ), .C(n6514), .D(\regX[22][0] ), 
        .Y(n6694) );
  NOR2X1 U4217 ( .A(n6704), .B(n6687), .Y(n6514) );
  INVX1 U4218 ( .A(n6518), .Y(n6619) );
  NAND3X1 U4219 ( .A(n6700), .B(n6698), .C(n6690), .Y(n6518) );
  INVX1 U4220 ( .A(n6705), .Y(n6690) );
  NOR2X1 U4221 ( .A(n6706), .B(n6707), .Y(n6678) );
  OAI21X1 U4222 ( .A(n3679), .B(n6622), .C(n6708), .Y(n6707) );
  AOI22X1 U4223 ( .A(n6589), .B(\regX[23][0] ), .C(n6502), .D(\regX[21][0] ), 
        .Y(n6708) );
  AND2X1 U4224 ( .A(n6709), .B(n6689), .Y(n6502) );
  NOR2X1 U4225 ( .A(n6710), .B(n6687), .Y(n6589) );
  INVX1 U4226 ( .A(n6497), .Y(n6622) );
  NOR2X1 U4227 ( .A(n6711), .B(n6687), .Y(n6497) );
  NAND2X1 U4228 ( .A(n6712), .B(n6713), .Y(n6706) );
  AOI22X1 U4229 ( .A(n6507), .B(\regX[19][0] ), .C(n6508), .D(\regX[13][0] ), 
        .Y(n6713) );
  AND2X1 U4230 ( .A(n6689), .B(n6692), .Y(n6508) );
  INVX1 U4231 ( .A(n6711), .Y(n6692) );
  NAND3X1 U4232 ( .A(n7205), .B(n6714), .C(n6715), .Y(n6711) );
  AND2X1 U4233 ( .A(n6709), .B(n6685), .Y(n6507) );
  AOI22X1 U4234 ( .A(n6509), .B(\regX[20][0] ), .C(n6626), .D(\regX[18][0] ), 
        .Y(n6712) );
  INVX1 U4235 ( .A(n6505), .Y(n6626) );
  NAND2X1 U4236 ( .A(n6685), .B(n6716), .Y(n6505) );
  NOR2X1 U4237 ( .A(n6717), .B(n6718), .Y(n6685) );
  AND2X1 U4238 ( .A(n6689), .B(n6716), .Y(n6509) );
  NOR2X1 U4239 ( .A(n6719), .B(n6720), .Y(n6677) );
  OAI21X1 U4240 ( .A(n3477), .B(n6201), .C(n6721), .Y(n6720) );
  AOI22X1 U4241 ( .A(n6494), .B(\regX[24][0] ), .C(n6630), .D(\regX[17][0] ), 
        .Y(n6721) );
  INVX1 U4242 ( .A(n6491), .Y(n6630) );
  NAND2X1 U4243 ( .A(n6709), .B(n6698), .Y(n6491) );
  INVX1 U4244 ( .A(n6710), .Y(n6709) );
  NAND3X1 U4245 ( .A(n7205), .B(n6722), .C(n6715), .Y(n6710) );
  INVX1 U4246 ( .A(n6723), .Y(n6494) );
  NAND3X1 U4247 ( .A(n6722), .B(n6714), .C(n7205), .Y(n6723) );
  OAI21X1 U4248 ( .A(n3666), .B(n6583), .C(n6724), .Y(n6719) );
  AOI22X1 U4249 ( .A(n6498), .B(N1735), .C(n6632), .D(N1433), .Y(n6724) );
  INVX1 U4250 ( .A(n6495), .Y(n6632) );
  NAND2X1 U4251 ( .A(n6689), .B(n6693), .Y(n6495) );
  INVX1 U4252 ( .A(n6688), .Y(n6693) );
  NAND3X1 U4253 ( .A(n6700), .B(n6701), .C(n6725), .Y(n6688) );
  NOR2X1 U4254 ( .A(n6715), .B(n6480), .Y(n6725) );
  AND2X1 U4255 ( .A(n6718), .B(n6717), .Y(n6689) );
  NOR2X1 U4256 ( .A(n6705), .B(n6687), .Y(n6498) );
  NAND2X1 U4257 ( .A(n6726), .B(n6718), .Y(n6687) );
  NAND3X1 U4258 ( .A(n6714), .B(n6703), .C(n7205), .Y(n6705) );
  NAND3X1 U4259 ( .A(n6701), .B(n6698), .C(n6716), .Y(n6583) );
  INVX1 U4260 ( .A(n6704), .Y(n6716) );
  NAND3X1 U4261 ( .A(n6722), .B(n6703), .C(n7205), .Y(n6704) );
  INVX1 U4262 ( .A(n6700), .Y(n6722) );
  XOR2X1 U4263 ( .A(n6727), .B(n6728), .Y(n6700) );
  XNOR2X1 U4264 ( .A(n6729), .B(n6730), .Y(n6727) );
  OAI21X1 U4265 ( .A(n6731), .B(n6732), .C(n6733), .Y(n6730) );
  OAI21X1 U4266 ( .A(n6734), .B(n6735), .C(n6728), .Y(n6733) );
  INVX1 U4267 ( .A(n6735), .Y(n6732) );
  OAI21X1 U4268 ( .A(n6736), .B(n6737), .C(n6738), .Y(n6729) );
  OAI21X1 U4269 ( .A(n6739), .B(n6740), .C(n6464), .Y(n6738) );
  NOR2X1 U4270 ( .A(n6741), .B(n6480), .Y(n6464) );
  NAND2X1 U4271 ( .A(n6742), .B(n6741), .Y(n6737) );
  INVX1 U4272 ( .A(N3343), .Y(n6741) );
  NOR2X1 U4273 ( .A(n6718), .B(n6726), .Y(n6698) );
  INVX1 U4274 ( .A(\regX[16][0] ), .Y(n3666) );
  NOR2X1 U4275 ( .A(n3477), .B(n4083), .Y(\U3/U118/Z_9 ) );
  INVX1 U4276 ( .A(fGy[9]), .Y(n4083) );
  NOR2X1 U4277 ( .A(n3477), .B(n4081), .Y(\U3/U118/Z_8 ) );
  INVX1 U4278 ( .A(fGy[8]), .Y(n4081) );
  OAI21X1 U4279 ( .A(n6743), .B(n5827), .C(n3529), .Y(\U3/U118/Z_7 ) );
  NAND2X1 U4280 ( .A(fGy[7]), .B(n3467), .Y(n3529) );
  NOR2X1 U4281 ( .A(n6744), .B(n6745), .Y(n6743) );
  NAND2X1 U4282 ( .A(n6746), .B(n6747), .Y(n6745) );
  NOR2X1 U4283 ( .A(n6748), .B(n6749), .Y(n6747) );
  OAI21X1 U4284 ( .A(n3849), .B(n6750), .C(n6751), .Y(n6749) );
  AOI22X1 U4285 ( .A(n6752), .B(\regX[11][7] ), .C(n6753), .D(\regX[7][7] ), 
        .Y(n6751) );
  OAI21X1 U4286 ( .A(n3922), .B(n6754), .C(n6755), .Y(n6748) );
  AOI22X1 U4287 ( .A(n6756), .B(N1622), .C(n6757), .D(\regX[23][7] ), .Y(n6755) );
  INVX1 U4288 ( .A(\regX[1][7] ), .Y(n3922) );
  NOR2X1 U4289 ( .A(n6758), .B(n6759), .Y(n6746) );
  OAI21X1 U4290 ( .A(n3813), .B(n6760), .C(n6761), .Y(n6759) );
  AOI22X1 U4291 ( .A(n6762), .B(\regX[5][7] ), .C(n6763), .D(\regX[0][7] ), 
        .Y(n6761) );
  INVX1 U4292 ( .A(\regX[9][7] ), .Y(n3813) );
  OAI21X1 U4293 ( .A(n3911), .B(n6764), .C(n6765), .Y(n6758) );
  AOI22X1 U4294 ( .A(n6766), .B(\regX[13][7] ), .C(n6767), .D(N1440), .Y(n6765) );
  NAND3X1 U4295 ( .A(n6768), .B(n6769), .C(n6770), .Y(n6744) );
  NOR2X1 U4296 ( .A(n6771), .B(n6772), .Y(n6770) );
  OAI21X1 U4297 ( .A(n3825), .B(n6773), .C(n6774), .Y(n6772) );
  AOI22X1 U4298 ( .A(n6775), .B(N1684), .C(n6776), .D(\regX[17][7] ), .Y(n6774) );
  INVX1 U4299 ( .A(\regX[8][7] ), .Y(n3825) );
  OAI21X1 U4300 ( .A(n3753), .B(n6777), .C(n6778), .Y(n6771) );
  AOI22X1 U4301 ( .A(n6779), .B(N1742), .C(n6780), .D(\regX[19][7] ), .Y(n6778) );
  INVX1 U4302 ( .A(\regX[15][7] ), .Y(n3753) );
  NOR2X1 U4303 ( .A(n6781), .B(n6782), .Y(n6769) );
  OAI22X1 U4304 ( .A(n3899), .B(n6783), .C(n3608), .D(n6784), .Y(n6782) );
  INVX1 U4305 ( .A(\regX[22][7] ), .Y(n3608) );
  INVX1 U4306 ( .A(\regX[3][7] ), .Y(n3899) );
  OAI22X1 U4307 ( .A(n3630), .B(n6785), .C(n3575), .D(n6786), .Y(n6781) );
  INVX1 U4308 ( .A(\regX[24][7] ), .Y(n3575) );
  INVX1 U4309 ( .A(\regX[20][7] ), .Y(n3630) );
  AOI21X1 U4310 ( .A(n6787), .B(\regX[16][7] ), .C(n6788), .Y(n6768) );
  OAI22X1 U4311 ( .A(n3651), .B(n6789), .C(n3619), .D(n6790), .Y(n6788) );
  INVX1 U4312 ( .A(\regX[21][7] ), .Y(n3619) );
  OAI21X1 U4313 ( .A(n6791), .B(n5827), .C(n3530), .Y(\U3/U118/Z_6 ) );
  NAND2X1 U4314 ( .A(fGy[6]), .B(n3467), .Y(n3530) );
  NOR2X1 U4315 ( .A(n6792), .B(n6793), .Y(n6791) );
  NAND2X1 U4316 ( .A(n6794), .B(n6795), .Y(n6793) );
  NOR2X1 U4317 ( .A(n6796), .B(n6797), .Y(n6795) );
  OAI21X1 U4318 ( .A(n3848), .B(n6750), .C(n6798), .Y(n6797) );
  AOI22X1 U4319 ( .A(n6752), .B(\regX[11][6] ), .C(n6753), .D(\regX[7][6] ), 
        .Y(n6798) );
  OAI21X1 U4320 ( .A(n3921), .B(n6754), .C(n6799), .Y(n6796) );
  AOI22X1 U4321 ( .A(n6756), .B(N1621), .C(n6757), .D(\regX[23][6] ), .Y(n6799) );
  INVX1 U4322 ( .A(\regX[1][6] ), .Y(n3921) );
  NOR2X1 U4323 ( .A(n6800), .B(n6801), .Y(n6794) );
  OAI21X1 U4324 ( .A(n3812), .B(n6760), .C(n6802), .Y(n6801) );
  AOI22X1 U4325 ( .A(n6762), .B(\regX[5][6] ), .C(n6763), .D(\regX[0][6] ), 
        .Y(n6802) );
  INVX1 U4326 ( .A(\regX[9][6] ), .Y(n3812) );
  OAI21X1 U4327 ( .A(n3910), .B(n6764), .C(n6803), .Y(n6800) );
  AOI22X1 U4328 ( .A(n6766), .B(\regX[13][6] ), .C(n6767), .D(N1439), .Y(n6803) );
  NAND3X1 U4329 ( .A(n6804), .B(n6805), .C(n6806), .Y(n6792) );
  NOR2X1 U4330 ( .A(n6807), .B(n6808), .Y(n6806) );
  OAI21X1 U4331 ( .A(n3824), .B(n6773), .C(n6809), .Y(n6808) );
  AOI22X1 U4332 ( .A(n6775), .B(N1683), .C(n6776), .D(\regX[17][6] ), .Y(n6809) );
  INVX1 U4333 ( .A(\regX[8][6] ), .Y(n3824) );
  OAI21X1 U4334 ( .A(n3752), .B(n6777), .C(n6810), .Y(n6807) );
  AOI22X1 U4335 ( .A(n6779), .B(N1741), .C(n6780), .D(\regX[19][6] ), .Y(n6810) );
  INVX1 U4336 ( .A(\regX[15][6] ), .Y(n3752) );
  NOR2X1 U4337 ( .A(n6811), .B(n6812), .Y(n6805) );
  OAI22X1 U4338 ( .A(n3898), .B(n6783), .C(n3607), .D(n6784), .Y(n6812) );
  INVX1 U4339 ( .A(\regX[22][6] ), .Y(n3607) );
  INVX1 U4340 ( .A(\regX[3][6] ), .Y(n3898) );
  OAI22X1 U4341 ( .A(n3629), .B(n6785), .C(n3573), .D(n6786), .Y(n6811) );
  INVX1 U4342 ( .A(\regX[24][6] ), .Y(n3573) );
  INVX1 U4343 ( .A(\regX[20][6] ), .Y(n3629) );
  AOI21X1 U4344 ( .A(n6787), .B(\regX[16][6] ), .C(n6813), .Y(n6804) );
  OAI22X1 U4345 ( .A(n3650), .B(n6789), .C(n3618), .D(n6790), .Y(n6813) );
  INVX1 U4346 ( .A(\regX[21][6] ), .Y(n3618) );
  OAI21X1 U4347 ( .A(n6814), .B(n5827), .C(n3531), .Y(\U3/U118/Z_5 ) );
  NAND2X1 U4348 ( .A(fGy[5]), .B(n3467), .Y(n3531) );
  NOR2X1 U4349 ( .A(n6815), .B(n6816), .Y(n6814) );
  NAND2X1 U4350 ( .A(n6817), .B(n6818), .Y(n6816) );
  NOR2X1 U4351 ( .A(n6819), .B(n6820), .Y(n6818) );
  OAI21X1 U4352 ( .A(n3847), .B(n6750), .C(n6821), .Y(n6820) );
  AOI22X1 U4353 ( .A(n6752), .B(\regX[11][5] ), .C(n6753), .D(\regX[7][5] ), 
        .Y(n6821) );
  INVX1 U4354 ( .A(\regX[6][5] ), .Y(n3847) );
  OAI21X1 U4355 ( .A(n3920), .B(n6754), .C(n6822), .Y(n6819) );
  AOI22X1 U4356 ( .A(n6756), .B(N1620), .C(n6757), .D(\regX[23][5] ), .Y(n6822) );
  INVX1 U4357 ( .A(\regX[1][5] ), .Y(n3920) );
  NOR2X1 U4358 ( .A(n6823), .B(n6824), .Y(n6817) );
  OAI21X1 U4359 ( .A(n3811), .B(n6760), .C(n6825), .Y(n6824) );
  AOI22X1 U4360 ( .A(n6762), .B(\regX[5][5] ), .C(n6763), .D(\regX[0][5] ), 
        .Y(n6825) );
  INVX1 U4361 ( .A(\regX[9][5] ), .Y(n3811) );
  OAI21X1 U4362 ( .A(n3909), .B(n6764), .C(n6826), .Y(n6823) );
  AOI22X1 U4363 ( .A(n6766), .B(\regX[13][5] ), .C(n6767), .D(N1438), .Y(n6826) );
  NAND3X1 U4364 ( .A(n6827), .B(n6828), .C(n6829), .Y(n6815) );
  NOR2X1 U4365 ( .A(n6830), .B(n6831), .Y(n6829) );
  OAI21X1 U4366 ( .A(n3823), .B(n6773), .C(n6832), .Y(n6831) );
  AOI22X1 U4367 ( .A(n6775), .B(N1682), .C(n6776), .D(\regX[17][5] ), .Y(n6832) );
  INVX1 U4368 ( .A(\regX[8][5] ), .Y(n3823) );
  OAI21X1 U4369 ( .A(n3751), .B(n6777), .C(n6833), .Y(n6830) );
  AOI22X1 U4370 ( .A(n6779), .B(N1740), .C(n6780), .D(\regX[19][5] ), .Y(n6833) );
  INVX1 U4371 ( .A(\regX[15][5] ), .Y(n3751) );
  NOR2X1 U4372 ( .A(n6834), .B(n6835), .Y(n6828) );
  OAI22X1 U4373 ( .A(n3897), .B(n6783), .C(n3606), .D(n6784), .Y(n6835) );
  INVX1 U4374 ( .A(\regX[22][5] ), .Y(n3606) );
  INVX1 U4375 ( .A(\regX[3][5] ), .Y(n3897) );
  OAI22X1 U4376 ( .A(n3628), .B(n6785), .C(n3571), .D(n6786), .Y(n6834) );
  INVX1 U4377 ( .A(\regX[24][5] ), .Y(n3571) );
  INVX1 U4378 ( .A(\regX[20][5] ), .Y(n3628) );
  AOI21X1 U4379 ( .A(n6787), .B(\regX[16][5] ), .C(n6836), .Y(n6827) );
  OAI22X1 U4380 ( .A(n3649), .B(n6789), .C(n3617), .D(n6790), .Y(n6836) );
  INVX1 U4381 ( .A(\regX[21][5] ), .Y(n3617) );
  OAI21X1 U4382 ( .A(n6837), .B(n5827), .C(n3532), .Y(\U3/U118/Z_4 ) );
  NAND2X1 U4383 ( .A(fGy[4]), .B(n3467), .Y(n3532) );
  NOR2X1 U4384 ( .A(n6838), .B(n6839), .Y(n6837) );
  NAND2X1 U4385 ( .A(n6840), .B(n6841), .Y(n6839) );
  NOR2X1 U4386 ( .A(n6842), .B(n6843), .Y(n6841) );
  OAI21X1 U4387 ( .A(n3846), .B(n6750), .C(n6844), .Y(n6843) );
  AOI22X1 U4388 ( .A(n6752), .B(\regX[11][4] ), .C(n6753), .D(\regX[7][4] ), 
        .Y(n6844) );
  OAI21X1 U4389 ( .A(n3919), .B(n6754), .C(n6845), .Y(n6842) );
  AOI22X1 U4390 ( .A(n6756), .B(N1619), .C(n6757), .D(\regX[23][4] ), .Y(n6845) );
  INVX1 U4391 ( .A(\regX[1][4] ), .Y(n3919) );
  NOR2X1 U4392 ( .A(n6846), .B(n6847), .Y(n6840) );
  OAI21X1 U4393 ( .A(n3810), .B(n6760), .C(n6848), .Y(n6847) );
  AOI22X1 U4394 ( .A(n6762), .B(\regX[5][4] ), .C(n6763), .D(\regX[0][4] ), 
        .Y(n6848) );
  INVX1 U4395 ( .A(\regX[9][4] ), .Y(n3810) );
  OAI21X1 U4396 ( .A(n3908), .B(n6764), .C(n6849), .Y(n6846) );
  AOI22X1 U4397 ( .A(n6766), .B(\regX[13][4] ), .C(n6767), .D(N1437), .Y(n6849) );
  NAND3X1 U4398 ( .A(n6850), .B(n6851), .C(n6852), .Y(n6838) );
  NOR2X1 U4399 ( .A(n6853), .B(n6854), .Y(n6852) );
  OAI21X1 U4400 ( .A(n3822), .B(n6773), .C(n6855), .Y(n6854) );
  AOI22X1 U4401 ( .A(n6775), .B(N1681), .C(n6776), .D(\regX[17][4] ), .Y(n6855) );
  INVX1 U4402 ( .A(\regX[8][4] ), .Y(n3822) );
  OAI21X1 U4403 ( .A(n3750), .B(n6777), .C(n6856), .Y(n6853) );
  AOI22X1 U4404 ( .A(n6779), .B(N1739), .C(n6780), .D(\regX[19][4] ), .Y(n6856) );
  INVX1 U4405 ( .A(\regX[15][4] ), .Y(n3750) );
  NOR2X1 U4406 ( .A(n6857), .B(n6858), .Y(n6851) );
  OAI22X1 U4407 ( .A(n3896), .B(n6783), .C(n3605), .D(n6784), .Y(n6858) );
  INVX1 U4408 ( .A(\regX[22][4] ), .Y(n3605) );
  INVX1 U4409 ( .A(\regX[3][4] ), .Y(n3896) );
  OAI22X1 U4410 ( .A(n3627), .B(n6785), .C(n3569), .D(n6786), .Y(n6857) );
  INVX1 U4411 ( .A(\regX[24][4] ), .Y(n3569) );
  INVX1 U4412 ( .A(\regX[20][4] ), .Y(n3627) );
  AOI21X1 U4413 ( .A(n6787), .B(\regX[16][4] ), .C(n6859), .Y(n6850) );
  OAI22X1 U4414 ( .A(n3648), .B(n6789), .C(n3616), .D(n6790), .Y(n6859) );
  INVX1 U4415 ( .A(\regX[21][4] ), .Y(n3616) );
  AND2X1 U4416 ( .A(n3467), .B(fGy[31]), .Y(\U3/U118/Z_31 ) );
  NOR2X1 U4417 ( .A(n3477), .B(n4125), .Y(\U3/U118/Z_30 ) );
  INVX1 U4418 ( .A(fGy[30]), .Y(n4125) );
  OAI21X1 U4419 ( .A(n3477), .B(n6479), .C(n6860), .Y(\U3/U118/Z_3 ) );
  AOI21X1 U4420 ( .A(n7246), .B(n6861), .C(n7205), .Y(n6860) );
  NAND3X1 U4421 ( .A(n6862), .B(n6863), .C(n6864), .Y(n6861) );
  NOR2X1 U4422 ( .A(n6865), .B(n6866), .Y(n6864) );
  OR2X1 U4423 ( .A(n6867), .B(n6868), .Y(n6866) );
  OAI21X1 U4424 ( .A(n3821), .B(n6773), .C(n6869), .Y(n6868) );
  AOI22X1 U4425 ( .A(n6775), .B(N1680), .C(n6776), .D(\regX[17][3] ), .Y(n6869) );
  INVX1 U4426 ( .A(\regX[8][3] ), .Y(n3821) );
  OAI21X1 U4427 ( .A(n3749), .B(n6777), .C(n6870), .Y(n6867) );
  AOI22X1 U4428 ( .A(n6779), .B(N1738), .C(n6780), .D(\regX[19][3] ), .Y(n6870) );
  INVX1 U4429 ( .A(\regX[15][3] ), .Y(n3749) );
  NAND3X1 U4430 ( .A(n6871), .B(n6872), .C(n6873), .Y(n6865) );
  AOI21X1 U4431 ( .A(n6787), .B(\regX[16][3] ), .C(n6874), .Y(n6873) );
  OAI22X1 U4432 ( .A(n3647), .B(n6789), .C(n3615), .D(n6790), .Y(n6874) );
  INVX1 U4433 ( .A(\regX[21][3] ), .Y(n3615) );
  AOI22X1 U4434 ( .A(n6875), .B(\regX[24][3] ), .C(n6876), .D(\regX[20][3] ), 
        .Y(n6872) );
  AOI22X1 U4435 ( .A(n6877), .B(\regX[22][3] ), .C(n6878), .D(\regX[3][3] ), 
        .Y(n6871) );
  NOR2X1 U4436 ( .A(n6879), .B(n6880), .Y(n6863) );
  OAI21X1 U4437 ( .A(n3845), .B(n6750), .C(n6881), .Y(n6880) );
  AOI22X1 U4438 ( .A(n6752), .B(\regX[11][3] ), .C(n6753), .D(\regX[7][3] ), 
        .Y(n6881) );
  OAI21X1 U4439 ( .A(n3918), .B(n6754), .C(n6882), .Y(n6879) );
  AOI22X1 U4440 ( .A(n6756), .B(N1618), .C(n6757), .D(\regX[23][3] ), .Y(n6882) );
  INVX1 U4441 ( .A(\regX[1][3] ), .Y(n3918) );
  NOR2X1 U4442 ( .A(n6883), .B(n6884), .Y(n6862) );
  OAI21X1 U4443 ( .A(n3809), .B(n6760), .C(n6885), .Y(n6884) );
  AOI22X1 U4444 ( .A(n6762), .B(\regX[5][3] ), .C(n6763), .D(\regX[0][3] ), 
        .Y(n6885) );
  INVX1 U4445 ( .A(\regX[9][3] ), .Y(n3809) );
  OAI21X1 U4446 ( .A(n3907), .B(n6764), .C(n6886), .Y(n6883) );
  AOI22X1 U4447 ( .A(n6766), .B(\regX[13][3] ), .C(n6767), .D(N1436), .Y(n6886) );
  NOR2X1 U4448 ( .A(n3477), .B(n4123), .Y(\U3/U118/Z_29 ) );
  INVX1 U4449 ( .A(fGy[29]), .Y(n4123) );
  NOR2X1 U4450 ( .A(n3477), .B(n4121), .Y(\U3/U118/Z_28 ) );
  INVX1 U4451 ( .A(fGy[28]), .Y(n4121) );
  NOR2X1 U4452 ( .A(n3477), .B(n4119), .Y(\U3/U118/Z_27 ) );
  INVX1 U4453 ( .A(fGy[27]), .Y(n4119) );
  NOR2X1 U4454 ( .A(n3477), .B(n4117), .Y(\U3/U118/Z_26 ) );
  INVX1 U4455 ( .A(fGy[26]), .Y(n4117) );
  NOR2X1 U4456 ( .A(n3477), .B(n4115), .Y(\U3/U118/Z_25 ) );
  INVX1 U4457 ( .A(fGy[25]), .Y(n4115) );
  NOR2X1 U4458 ( .A(n3477), .B(n4113), .Y(\U3/U118/Z_24 ) );
  INVX1 U4459 ( .A(fGy[24]), .Y(n4113) );
  NOR2X1 U4460 ( .A(n3477), .B(n4111), .Y(\U3/U118/Z_23 ) );
  INVX1 U4461 ( .A(fGy[23]), .Y(n4111) );
  NOR2X1 U4462 ( .A(n3477), .B(n4109), .Y(\U3/U118/Z_22 ) );
  INVX1 U4463 ( .A(fGy[22]), .Y(n4109) );
  NOR2X1 U4464 ( .A(n3477), .B(n4107), .Y(\U3/U118/Z_21 ) );
  INVX1 U4465 ( .A(fGy[21]), .Y(n4107) );
  NOR2X1 U4466 ( .A(n3477), .B(n4105), .Y(\U3/U118/Z_20 ) );
  INVX1 U4467 ( .A(fGy[20]), .Y(n4105) );
  NAND3X1 U4468 ( .A(n6480), .B(n3533), .C(n6887), .Y(\U3/U118/Z_2 ) );
  OAI21X1 U4469 ( .A(n6888), .B(n6889), .C(n7246), .Y(n6887) );
  NAND2X1 U4470 ( .A(n6890), .B(n6891), .Y(n6889) );
  NOR2X1 U4471 ( .A(n6892), .B(n6893), .Y(n6891) );
  OAI21X1 U4472 ( .A(n3844), .B(n6750), .C(n6894), .Y(n6893) );
  AOI22X1 U4473 ( .A(n6752), .B(\regX[11][2] ), .C(n6753), .D(\regX[7][2] ), 
        .Y(n6894) );
  OAI21X1 U4474 ( .A(n3917), .B(n6754), .C(n6895), .Y(n6892) );
  AOI22X1 U4475 ( .A(n6756), .B(N1617), .C(n6757), .D(\regX[23][2] ), .Y(n6895) );
  INVX1 U4476 ( .A(\regX[1][2] ), .Y(n3917) );
  NOR2X1 U4477 ( .A(n6896), .B(n6897), .Y(n6890) );
  OAI21X1 U4478 ( .A(n3808), .B(n6760), .C(n6898), .Y(n6897) );
  AOI22X1 U4479 ( .A(n6762), .B(\regX[5][2] ), .C(n6763), .D(\regX[0][2] ), 
        .Y(n6898) );
  INVX1 U4480 ( .A(\regX[9][2] ), .Y(n3808) );
  OAI21X1 U4481 ( .A(n3906), .B(n6764), .C(n6899), .Y(n6896) );
  AOI22X1 U4482 ( .A(n6766), .B(\regX[13][2] ), .C(n6767), .D(N1435), .Y(n6899) );
  NAND3X1 U4483 ( .A(n6900), .B(n6901), .C(n6902), .Y(n6888) );
  NOR2X1 U4484 ( .A(n6903), .B(n6904), .Y(n6902) );
  OAI21X1 U4485 ( .A(n3820), .B(n6773), .C(n6905), .Y(n6904) );
  AOI22X1 U4486 ( .A(n6775), .B(N1679), .C(n6776), .D(\regX[17][2] ), .Y(n6905) );
  INVX1 U4487 ( .A(\regX[8][2] ), .Y(n3820) );
  OAI21X1 U4488 ( .A(n3740), .B(n6777), .C(n6906), .Y(n6903) );
  AOI22X1 U4489 ( .A(n6779), .B(N1737), .C(n6780), .D(\regX[19][2] ), .Y(n6906) );
  INVX1 U4490 ( .A(\regX[15][2] ), .Y(n3740) );
  NOR2X1 U4491 ( .A(n6907), .B(n6908), .Y(n6901) );
  OAI22X1 U4492 ( .A(n3894), .B(n6783), .C(n3603), .D(n6784), .Y(n6908) );
  INVX1 U4493 ( .A(\regX[22][2] ), .Y(n3603) );
  INVX1 U4494 ( .A(\regX[3][2] ), .Y(n3894) );
  OAI22X1 U4495 ( .A(n3625), .B(n6785), .C(n3565), .D(n6786), .Y(n6907) );
  INVX1 U4496 ( .A(\regX[24][2] ), .Y(n3565) );
  INVX1 U4497 ( .A(\regX[20][2] ), .Y(n3625) );
  AOI21X1 U4498 ( .A(n6787), .B(\regX[16][2] ), .C(n6909), .Y(n6900) );
  OAI22X1 U4499 ( .A(n3646), .B(n6789), .C(n3614), .D(n6790), .Y(n6909) );
  INVX1 U4500 ( .A(\regX[21][2] ), .Y(n3614) );
  NAND2X1 U4501 ( .A(fGy[2]), .B(n3467), .Y(n3533) );
  NOR2X1 U4502 ( .A(n3477), .B(n4103), .Y(\U3/U118/Z_19 ) );
  INVX1 U4503 ( .A(fGy[19]), .Y(n4103) );
  NOR2X1 U4504 ( .A(n3477), .B(n4101), .Y(\U3/U118/Z_18 ) );
  INVX1 U4505 ( .A(fGy[18]), .Y(n4101) );
  NOR2X1 U4506 ( .A(n3477), .B(n4099), .Y(\U3/U118/Z_17 ) );
  INVX1 U4507 ( .A(fGy[17]), .Y(n4099) );
  NOR2X1 U4508 ( .A(n3477), .B(n4097), .Y(\U3/U118/Z_16 ) );
  INVX1 U4509 ( .A(fGy[16]), .Y(n4097) );
  NOR2X1 U4510 ( .A(n3477), .B(n4095), .Y(\U3/U118/Z_15 ) );
  INVX1 U4511 ( .A(fGy[15]), .Y(n4095) );
  NOR2X1 U4512 ( .A(n3477), .B(n4093), .Y(\U3/U118/Z_14 ) );
  INVX1 U4513 ( .A(fGy[14]), .Y(n4093) );
  NOR2X1 U4514 ( .A(n3477), .B(n4091), .Y(\U3/U118/Z_13 ) );
  INVX1 U4515 ( .A(fGy[13]), .Y(n4091) );
  NOR2X1 U4516 ( .A(n3477), .B(n4089), .Y(\U3/U118/Z_12 ) );
  INVX1 U4517 ( .A(fGy[12]), .Y(n4089) );
  NOR2X1 U4518 ( .A(n3477), .B(n4087), .Y(\U3/U118/Z_11 ) );
  INVX1 U4519 ( .A(fGy[11]), .Y(n4087) );
  NOR2X1 U4520 ( .A(n3477), .B(n4085), .Y(\U3/U118/Z_10 ) );
  INVX1 U4521 ( .A(fGy[10]), .Y(n4085) );
  OAI21X1 U4522 ( .A(n3477), .B(n6482), .C(n6910), .Y(\U3/U118/Z_1 ) );
  AOI21X1 U4523 ( .A(n7246), .B(n6911), .C(n7205), .Y(n6910) );
  NAND3X1 U4524 ( .A(n6912), .B(n6913), .C(n6914), .Y(n6911) );
  NOR2X1 U4525 ( .A(n6915), .B(n6916), .Y(n6914) );
  OR2X1 U4526 ( .A(n6917), .B(n6918), .Y(n6916) );
  OAI21X1 U4527 ( .A(n3819), .B(n6773), .C(n6919), .Y(n6918) );
  AOI22X1 U4528 ( .A(n6775), .B(N1678), .C(n6776), .D(\regX[17][1] ), .Y(n6919) );
  INVX1 U4529 ( .A(\regX[8][1] ), .Y(n3819) );
  OAI21X1 U4530 ( .A(n3681), .B(n6777), .C(n6920), .Y(n6917) );
  AOI22X1 U4531 ( .A(n6779), .B(N1736), .C(n6780), .D(\regX[19][1] ), .Y(n6920) );
  INVX1 U4532 ( .A(\regX[15][1] ), .Y(n3681) );
  NAND3X1 U4533 ( .A(n6921), .B(n6922), .C(n6923), .Y(n6915) );
  AOI21X1 U4534 ( .A(n6787), .B(\regX[16][1] ), .C(n6924), .Y(n6923) );
  OAI22X1 U4535 ( .A(n3645), .B(n6789), .C(n3613), .D(n6790), .Y(n6924) );
  INVX1 U4536 ( .A(\regX[21][1] ), .Y(n3613) );
  AOI22X1 U4537 ( .A(n6875), .B(\regX[24][1] ), .C(n6876), .D(\regX[20][1] ), 
        .Y(n6922) );
  INVX1 U4538 ( .A(n6785), .Y(n6876) );
  AOI22X1 U4539 ( .A(n6877), .B(\regX[22][1] ), .C(n6878), .D(\regX[3][1] ), 
        .Y(n6921) );
  INVX1 U4540 ( .A(n6783), .Y(n6878) );
  INVX1 U4541 ( .A(n6784), .Y(n6877) );
  NOR2X1 U4542 ( .A(n6925), .B(n6926), .Y(n6913) );
  OAI21X1 U4543 ( .A(n3843), .B(n6750), .C(n6927), .Y(n6926) );
  AOI22X1 U4544 ( .A(n6752), .B(\regX[11][1] ), .C(n6753), .D(\regX[7][1] ), 
        .Y(n6927) );
  OAI21X1 U4545 ( .A(n3916), .B(n6754), .C(n6928), .Y(n6925) );
  AOI22X1 U4546 ( .A(n6756), .B(N1616), .C(n6757), .D(\regX[23][1] ), .Y(n6928) );
  INVX1 U4547 ( .A(\regX[1][1] ), .Y(n3916) );
  NOR2X1 U4548 ( .A(n6929), .B(n6930), .Y(n6912) );
  OAI21X1 U4549 ( .A(n3807), .B(n6760), .C(n6931), .Y(n6930) );
  AOI22X1 U4550 ( .A(n6762), .B(\regX[5][1] ), .C(n6763), .D(\regX[0][1] ), 
        .Y(n6931) );
  INVX1 U4551 ( .A(\regX[9][1] ), .Y(n3807) );
  OAI21X1 U4552 ( .A(n3905), .B(n6764), .C(n6932), .Y(n6929) );
  AOI22X1 U4553 ( .A(n6766), .B(\regX[13][1] ), .C(n6767), .D(N1434), .Y(n6932) );
  NAND3X1 U4554 ( .A(n6480), .B(n3534), .C(n6933), .Y(\U3/U118/Z_0 ) );
  OAI21X1 U4555 ( .A(n6934), .B(n6935), .C(n7246), .Y(n6933) );
  NAND2X1 U4556 ( .A(n6936), .B(n6937), .Y(n6935) );
  NOR2X1 U4557 ( .A(n6938), .B(n6939), .Y(n6937) );
  OAI21X1 U4558 ( .A(n3841), .B(n6750), .C(n6940), .Y(n6939) );
  AOI22X1 U4559 ( .A(n6752), .B(\regX[11][0] ), .C(n6753), .D(\regX[7][0] ), 
        .Y(n6940) );
  AND2X1 U4560 ( .A(n6941), .B(n6942), .Y(n6753) );
  AND2X1 U4561 ( .A(n6943), .B(n6944), .Y(n6752) );
  NAND2X1 U4562 ( .A(n6945), .B(n6942), .Y(n6750) );
  OAI21X1 U4563 ( .A(n3914), .B(n6754), .C(n6946), .Y(n6938) );
  AOI22X1 U4564 ( .A(n6756), .B(N1615), .C(n6757), .D(\regX[23][0] ), .Y(n6946) );
  AND2X1 U4565 ( .A(n6947), .B(n6942), .Y(n6757) );
  AND2X1 U4566 ( .A(n6948), .B(n6944), .Y(n6756) );
  NAND2X1 U4567 ( .A(n6949), .B(n6941), .Y(n6754) );
  INVX1 U4568 ( .A(\regX[1][0] ), .Y(n3914) );
  NOR2X1 U4569 ( .A(n6950), .B(n6951), .Y(n6936) );
  OAI21X1 U4570 ( .A(n3805), .B(n6760), .C(n6952), .Y(n6951) );
  AOI22X1 U4571 ( .A(n6762), .B(\regX[5][0] ), .C(n6763), .D(\regX[0][0] ), 
        .Y(n6952) );
  AND2X1 U4572 ( .A(n6945), .B(n6949), .Y(n6763) );
  AND2X1 U4573 ( .A(n6941), .B(n6953), .Y(n6762) );
  NAND2X1 U4574 ( .A(n6943), .B(n6949), .Y(n6760) );
  INVX1 U4575 ( .A(\regX[9][0] ), .Y(n3805) );
  OAI21X1 U4576 ( .A(n3903), .B(n6764), .C(n6954), .Y(n6950) );
  AOI22X1 U4577 ( .A(n6766), .B(\regX[13][0] ), .C(n6767), .D(N1433), .Y(n6954) );
  AND2X1 U4578 ( .A(n6945), .B(n6953), .Y(n6767) );
  AND2X1 U4579 ( .A(n6943), .B(n6953), .Y(n6766) );
  NAND2X1 U4580 ( .A(n6945), .B(n6944), .Y(n6764) );
  INVX1 U4581 ( .A(n6955), .Y(n6945) );
  NAND3X1 U4582 ( .A(n6956), .B(n6957), .C(n6958), .Y(n6955) );
  INVX1 U4583 ( .A(N1375), .Y(n3903) );
  NAND3X1 U4584 ( .A(n6959), .B(n6960), .C(n6961), .Y(n6934) );
  NOR2X1 U4585 ( .A(n6962), .B(n6963), .Y(n6961) );
  OAI21X1 U4586 ( .A(n3817), .B(n6773), .C(n6964), .Y(n6963) );
  AOI22X1 U4587 ( .A(n6775), .B(N1677), .C(n6776), .D(\regX[17][0] ), .Y(n6964) );
  AND2X1 U4588 ( .A(n6949), .B(n6947), .Y(n6776) );
  AND2X1 U4589 ( .A(n6948), .B(n6953), .Y(n6775) );
  NAND3X1 U4590 ( .A(n6949), .B(n6958), .C(n6948), .Y(n6773) );
  INVX1 U4591 ( .A(\regX[8][0] ), .Y(n3817) );
  OAI21X1 U4592 ( .A(n3679), .B(n6777), .C(n6965), .Y(n6962) );
  AOI22X1 U4593 ( .A(n6779), .B(N1735), .C(n6780), .D(\regX[19][0] ), .Y(n6965) );
  AND2X1 U4594 ( .A(n6947), .B(n6944), .Y(n6780) );
  AND2X1 U4595 ( .A(n6948), .B(n6942), .Y(n6779) );
  NOR2X1 U4596 ( .A(n6956), .B(n6966), .Y(n6948) );
  NAND2X1 U4597 ( .A(n6943), .B(n6942), .Y(n6777) );
  NOR2X1 U4598 ( .A(n6957), .B(n6956), .Y(n6943) );
  INVX1 U4599 ( .A(\regX[15][0] ), .Y(n3679) );
  NOR2X1 U4600 ( .A(n6967), .B(n6968), .Y(n6960) );
  OAI22X1 U4601 ( .A(n3891), .B(n6783), .C(n3600), .D(n6784), .Y(n6968) );
  NAND2X1 U4602 ( .A(n6942), .B(n6969), .Y(n6784) );
  AND2X1 U4603 ( .A(n6970), .B(n6971), .Y(n6942) );
  INVX1 U4604 ( .A(\regX[22][0] ), .Y(n3600) );
  NAND2X1 U4605 ( .A(n6944), .B(n6941), .Y(n6783) );
  INVX1 U4606 ( .A(n6972), .Y(n6941) );
  NAND3X1 U4607 ( .A(n6958), .B(n6956), .C(n6966), .Y(n6972) );
  INVX1 U4608 ( .A(\regX[3][0] ), .Y(n3891) );
  OAI22X1 U4609 ( .A(n3622), .B(n6785), .C(n3560), .D(n6786), .Y(n6967) );
  INVX1 U4610 ( .A(n6875), .Y(n6786) );
  NOR2X1 U4611 ( .A(n6956), .B(n6958), .Y(n6875) );
  INVX1 U4612 ( .A(\regX[24][0] ), .Y(n3560) );
  NAND2X1 U4613 ( .A(n6953), .B(n6969), .Y(n6785) );
  INVX1 U4614 ( .A(\regX[20][0] ), .Y(n3622) );
  AOI21X1 U4615 ( .A(n6787), .B(\regX[16][0] ), .C(n6973), .Y(n6959) );
  OAI22X1 U4616 ( .A(n3643), .B(n6789), .C(n3611), .D(n6790), .Y(n6973) );
  NAND2X1 U4617 ( .A(n6947), .B(n6953), .Y(n6790) );
  AND2X1 U4618 ( .A(n6974), .B(n6971), .Y(n6953) );
  NOR2X1 U4619 ( .A(n6957), .B(n6958), .Y(n6947) );
  INVX1 U4620 ( .A(\regX[21][0] ), .Y(n3611) );
  NAND2X1 U4621 ( .A(n6944), .B(n6969), .Y(n6789) );
  NOR2X1 U4622 ( .A(n6971), .B(n6974), .Y(n6944) );
  INVX1 U4623 ( .A(n6970), .Y(n6974) );
  INVX1 U4624 ( .A(n6975), .Y(n6787) );
  NAND3X1 U4625 ( .A(n6969), .B(n6956), .C(n6949), .Y(n6975) );
  NOR2X1 U4626 ( .A(n6971), .B(n6970), .Y(n6949) );
  XOR2X1 U4627 ( .A(n6451), .B(n6976), .Y(n6970) );
  XOR2X1 U4628 ( .A(N3090), .B(n6977), .Y(n6976) );
  OAI21X1 U4629 ( .A(n6978), .B(n6979), .C(n6980), .Y(n6971) );
  OAI21X1 U4630 ( .A(N3092), .B(n6980), .C(n6981), .Y(n6956) );
  NOR2X1 U4631 ( .A(n6958), .B(n6966), .Y(n6969) );
  INVX1 U4632 ( .A(n6957), .Y(n6966) );
  OAI21X1 U4633 ( .A(N3089), .B(n6447), .C(n6982), .Y(n6957) );
  XNOR2X1 U4634 ( .A(n6983), .B(N3093), .Y(n6958) );
  NAND2X1 U4635 ( .A(n6444), .B(n6981), .Y(n6983) );
  NAND2X1 U4636 ( .A(N3092), .B(n6980), .Y(n6981) );
  NAND2X1 U4637 ( .A(n6978), .B(n6979), .Y(n6980) );
  INVX1 U4638 ( .A(N3091), .Y(n6979) );
  INVX1 U4639 ( .A(n6984), .Y(n6978) );
  OAI21X1 U4640 ( .A(n6454), .B(n6982), .C(n6985), .Y(n6984) );
  OAI21X1 U4641 ( .A(n6977), .B(n6451), .C(N3090), .Y(n6985) );
  INVX1 U4642 ( .A(n6982), .Y(n6977) );
  NAND2X1 U4643 ( .A(N3089), .B(n6447), .Y(n6982) );
  INVX1 U4644 ( .A(n6445), .Y(n6447) );
  XNOR2X1 U4645 ( .A(n6986), .B(n6987), .Y(n6445) );
  NOR2X1 U4646 ( .A(n6480), .B(n6068), .Y(n6987) );
  INVX1 U4647 ( .A(n6451), .Y(n6454) );
  XOR2X1 U4648 ( .A(n6460), .B(n6988), .Y(n6451) );
  XOR2X1 U4649 ( .A(n6989), .B(n6990), .Y(n6988) );
  NAND2X1 U4650 ( .A(n6076), .B(n5827), .Y(n6990) );
  XNOR2X1 U4651 ( .A(n6991), .B(n6476), .Y(n6444) );
  XOR2X1 U4652 ( .A(n6472), .B(n6471), .Y(n6991) );
  INVX1 U4653 ( .A(n6475), .Y(n6471) );
  OAI21X1 U4654 ( .A(n6478), .B(n6075), .C(n6992), .Y(n6475) );
  OAI21X1 U4655 ( .A(n6082), .B(n6993), .C(n6476), .Y(n6992) );
  INVX1 U4656 ( .A(n6075), .Y(n6082) );
  XOR2X1 U4657 ( .A(n6994), .B(n6995), .Y(n6075) );
  XOR2X1 U4658 ( .A(n6996), .B(n6997), .Y(n6994) );
  INVX1 U4659 ( .A(n6993), .Y(n6478) );
  OAI21X1 U4660 ( .A(n6460), .B(n6989), .C(n6998), .Y(n6993) );
  OAI22X1 U4661 ( .A(n7246), .B(n6081), .C(n6999), .D(n6476), .Y(n6998) );
  INVX1 U4662 ( .A(n6989), .Y(n6999) );
  INVX1 U4663 ( .A(n6076), .Y(n6081) );
  XOR2X1 U4664 ( .A(n7000), .B(n7001), .Y(n6076) );
  XOR2X1 U4665 ( .A(n7002), .B(n7003), .Y(n7001) );
  OAI21X1 U4666 ( .A(n6068), .B(n6986), .C(n7205), .Y(n6989) );
  XOR2X1 U4667 ( .A(n6480), .B(n7004), .Y(n6986) );
  OAI21X1 U4668 ( .A(n7005), .B(n7006), .C(n7000), .Y(n6068) );
  NAND2X1 U4669 ( .A(n6715), .B(n7246), .Y(n7006) );
  INVX1 U4670 ( .A(n6476), .Y(n6460) );
  XNOR2X1 U4671 ( .A(n6480), .B(dx[1]), .Y(n6476) );
  NAND2X1 U4672 ( .A(n6064), .B(n7205), .Y(n6472) );
  XOR2X1 U4673 ( .A(n7007), .B(n6469), .Y(n6064) );
  INVX1 U4674 ( .A(n6465), .Y(n6469) );
  OAI21X1 U4675 ( .A(n5827), .B(n7008), .C(n6736), .Y(n6465) );
  INVX1 U4676 ( .A(N3092), .Y(n7008) );
  XOR2X1 U4677 ( .A(n6468), .B(n6470), .Y(n7007) );
  OAI21X1 U4678 ( .A(n7009), .B(n6995), .C(n7010), .Y(n6470) );
  OAI21X1 U4679 ( .A(n6996), .B(n7011), .C(n6997), .Y(n7010) );
  AOI21X1 U4680 ( .A(n7246), .B(N3091), .C(n7012), .Y(n6997) );
  INVX1 U4681 ( .A(n7009), .Y(n6996) );
  INVX1 U4682 ( .A(n7011), .Y(n6995) );
  OAI21X1 U4683 ( .A(n7003), .B(n7013), .C(n7014), .Y(n7011) );
  OAI21X1 U4684 ( .A(n7002), .B(n7015), .C(n7000), .Y(n7014) );
  OAI21X1 U4685 ( .A(n5827), .B(n6703), .C(n7005), .Y(n7000) );
  INVX1 U4686 ( .A(n7016), .Y(n7005) );
  AOI22X1 U4687 ( .A(n7205), .B(N3359), .C(n7246), .D(N3089), .Y(n7016) );
  INVX1 U4688 ( .A(n6715), .Y(n6703) );
  XNOR2X1 U4689 ( .A(n7017), .B(n7018), .Y(n6715) );
  NOR2X1 U4690 ( .A(N3359), .B(n7246), .Y(n7018) );
  INVX1 U4691 ( .A(n7002), .Y(n7013) );
  AOI21X1 U4692 ( .A(n7246), .B(N3090), .C(n7019), .Y(n7002) );
  INVX1 U4693 ( .A(n7015), .Y(n7003) );
  NAND2X1 U4694 ( .A(n6717), .B(n6480), .Y(n7015) );
  INVX1 U4695 ( .A(n6726), .Y(n6717) );
  XOR2X1 U4696 ( .A(n7020), .B(n6728), .Y(n6726) );
  XNOR2X1 U4697 ( .A(n7021), .B(n7022), .Y(n7020) );
  NAND2X1 U4698 ( .A(N3340), .B(n5827), .Y(n7021) );
  NOR2X1 U4699 ( .A(n6718), .B(n7205), .Y(n7009) );
  XNOR2X1 U4700 ( .A(n7023), .B(n6728), .Y(n6718) );
  XOR2X1 U4701 ( .A(n7024), .B(n7025), .Y(n7023) );
  INVX1 U4702 ( .A(n6466), .Y(n6468) );
  NAND2X1 U4703 ( .A(n7246), .B(n6714), .Y(n6466) );
  INVX1 U4704 ( .A(n6701), .Y(n6714) );
  XOR2X1 U4705 ( .A(n7026), .B(n6728), .Y(n6701) );
  XOR2X1 U4706 ( .A(n6735), .B(n6731), .Y(n7026) );
  INVX1 U4707 ( .A(n6734), .Y(n6731) );
  OAI21X1 U4708 ( .A(n7027), .B(n7025), .C(n7028), .Y(n6734) );
  OAI21X1 U4709 ( .A(n7024), .B(n7029), .C(n6728), .Y(n7028) );
  INVX1 U4710 ( .A(n7029), .Y(n7025) );
  OAI21X1 U4711 ( .A(n7030), .B(n7031), .C(n7032), .Y(n7029) );
  NOR2X1 U4712 ( .A(n6739), .B(n7246), .Y(n7032) );
  INVX1 U4713 ( .A(n7024), .Y(n7027) );
  OAI21X1 U4714 ( .A(n7033), .B(n7022), .C(n7034), .Y(n7024) );
  INVX1 U4715 ( .A(n7035), .Y(n7034) );
  AOI22X1 U4716 ( .A(n5827), .B(N3340), .C(n7022), .D(n7033), .Y(n7035) );
  OAI21X1 U4717 ( .A(n7246), .B(N3359), .C(n7017), .Y(n7022) );
  XOR2X1 U4718 ( .A(n5827), .B(n7004), .Y(n7017) );
  INVX1 U4719 ( .A(n6728), .Y(n7033) );
  XNOR2X1 U4720 ( .A(n5827), .B(dx[1]), .Y(n6728) );
  OAI21X1 U4721 ( .A(n6736), .B(n6742), .C(n7036), .Y(n6735) );
  OAI21X1 U4722 ( .A(n7012), .B(n7019), .C(n6740), .Y(n7036) );
  INVX1 U4723 ( .A(N3342), .Y(n6740) );
  INVX1 U4724 ( .A(n7031), .Y(n7019) );
  NAND2X1 U4725 ( .A(N3340), .B(n7205), .Y(n7031) );
  NOR2X1 U4726 ( .A(n7030), .B(n6480), .Y(n7012) );
  INVX1 U4727 ( .A(N3341), .Y(n7030) );
  INVX1 U4728 ( .A(n6739), .Y(n6742) );
  NOR2X1 U4729 ( .A(N3340), .B(N3341), .Y(n6739) );
  NAND2X1 U4730 ( .A(N3342), .B(n7205), .Y(n6736) );
  NAND2X1 U4731 ( .A(fGy[0]), .B(n3467), .Y(n3534) );
  OAI21X1 U4732 ( .A(n3475), .B(n3651), .C(n7037), .Y(\U3/U110/Z_7 ) );
  INVX1 U4733 ( .A(\regX[18][7] ), .Y(n3651) );
  OAI21X1 U4734 ( .A(n3475), .B(n3650), .C(n7037), .Y(\U3/U110/Z_6 ) );
  INVX1 U4735 ( .A(\regX[18][6] ), .Y(n3650) );
  OAI21X1 U4736 ( .A(n3475), .B(n3649), .C(n7037), .Y(\U3/U110/Z_5 ) );
  INVX1 U4737 ( .A(\regX[18][5] ), .Y(n3649) );
  OAI21X1 U4738 ( .A(n3475), .B(n3648), .C(n7037), .Y(\U3/U110/Z_4 ) );
  INVX1 U4739 ( .A(\regX[18][4] ), .Y(n3648) );
  OAI21X1 U4740 ( .A(n3475), .B(n3647), .C(n7037), .Y(\U3/U110/Z_3 ) );
  INVX1 U4741 ( .A(\regX[18][3] ), .Y(n3647) );
  OAI21X1 U4742 ( .A(n3475), .B(n3646), .C(n7037), .Y(\U3/U110/Z_2 ) );
  INVX1 U4743 ( .A(\regX[18][2] ), .Y(n3646) );
  OAI21X1 U4744 ( .A(n3475), .B(n3645), .C(n7037), .Y(\U3/U110/Z_1 ) );
  NAND2X1 U4745 ( .A(dy[1]), .B(n7205), .Y(n7037) );
  INVX1 U4746 ( .A(\regX[18][1] ), .Y(n3645) );
  OAI22X1 U4747 ( .A(n6480), .B(n5825), .C(n3475), .D(n3643), .Y(\U3/U110/Z_0 ) );
  INVX1 U4748 ( .A(\regX[18][0] ), .Y(n3643) );
  INVX1 U4749 ( .A(dy[0]), .Y(n5825) );
  NAND2X1 U4750 ( .A(n6480), .B(n3475), .Y(\U3/U109/Z_2 ) );
  NAND3X1 U4751 ( .A(n4257), .B(n4250), .C(n5724), .Y(n5823) );
  NOR2X1 U4752 ( .A(OPMode[2]), .B(OPMode[1]), .Y(n5724) );
  NAND2X1 U4753 ( .A(n3540), .B(n3554), .Y(n3548) );
  OAI21X1 U4754 ( .A(n3477), .B(n6479), .C(n7038), .Y(\U3/U106/Z_3 ) );
  INVX1 U4755 ( .A(fGy[3]), .Y(n6479) );
  OAI21X1 U4756 ( .A(n3477), .B(n6482), .C(n7038), .Y(\U3/U106/Z_1 ) );
  INVX1 U4757 ( .A(fGy[1]), .Y(n6482) );
  OAI22X1 U4758 ( .A(n3845), .B(n7038), .C(n3477), .D(n6176), .Y(\U3/U105/Z_3 ) );
  INVX1 U4759 ( .A(N2749), .Y(n6176) );
  INVX1 U4760 ( .A(\regX[6][3] ), .Y(n3845) );
  OAI22X1 U4761 ( .A(n3844), .B(n7038), .C(n3477), .D(n6179), .Y(\U3/U105/Z_2 ) );
  INVX1 U4762 ( .A(N2748), .Y(n6179) );
  INVX1 U4763 ( .A(\regX[6][2] ), .Y(n3844) );
  OAI22X1 U4764 ( .A(n3843), .B(n7038), .C(n3477), .D(n6190), .Y(\U3/U105/Z_1 ) );
  INVX1 U4765 ( .A(N2747), .Y(n6190) );
  INVX1 U4766 ( .A(\regX[6][1] ), .Y(n3843) );
  OAI22X1 U4767 ( .A(n3841), .B(n7038), .C(n3477), .D(n6201), .Y(\U3/U105/Z_0 ) );
  INVX1 U4768 ( .A(N2746), .Y(n6201) );
  INVX1 U4769 ( .A(n4612), .Y(n7038) );
  INVX1 U4770 ( .A(\regX[6][0] ), .Y(n3841) );
  NOR2X1 U4771 ( .A(n5692), .B(n4619), .Y(\U3/U101/Z_6 ) );
  XOR2X1 U4772 ( .A(n7039), .B(n4412), .Y(n4619) );
  OAI21X1 U4773 ( .A(n5161), .B(n7040), .C(n7041), .Y(n4412) );
  XOR2X1 U4774 ( .A(n5161), .B(n7042), .Y(n7039) );
  NOR2X1 U4775 ( .A(n7043), .B(n7044), .Y(n7042) );
  INVX1 U4776 ( .A(n5810), .Y(n7043) );
  NOR2X1 U4777 ( .A(n4683), .B(n5692), .Y(\U3/U101/Z_3 ) );
  INVX1 U4778 ( .A(bCE), .Y(n5692) );
  XOR2X1 U4779 ( .A(n7044), .B(n5810), .Y(n4683) );
  NAND2X1 U4780 ( .A(n5165), .B(n5809), .Y(n5810) );
  XOR2X1 U4781 ( .A(n5172), .B(n5161), .Y(n5809) );
  OAI21X1 U4782 ( .A(n5161), .B(n7045), .C(n7041), .Y(n5172) );
  INVX1 U4783 ( .A(N3441), .Y(n7045) );
  MUX2X1 U4784 ( .B(n5175), .A(n7046), .S(n7202), .Y(n5165) );
  NAND2X1 U4785 ( .A(n5174), .B(n5175), .Y(n7046) );
  OAI21X1 U4786 ( .A(n5161), .B(n7047), .C(n7041), .Y(n5175) );
  INVX1 U4787 ( .A(N1389), .Y(n7047) );
  XNOR2X1 U4790 ( .A(n4685), .B(n7202), .Y(n7044) );
  OAI21X1 U4791 ( .A(n5161), .B(n7048), .C(n7041), .Y(n4685) );
  NAND2X1 U4792 ( .A(dx[1]), .B(n7204), .Y(n7041) );
  INVX1 U4793 ( .A(n3943), .Y(n7204) );
  INVX1 U4794 ( .A(n7049), .Y(\U3/U101/Z_0 ) );
  MUX2X1 U4795 ( .B(dAddrRegCol[0]), .A(n5174), .S(bCE), .Y(n7049) );
  OAI21X1 U4796 ( .A(n3943), .B(n7004), .C(n7050), .Y(n5174) );
  NAND2X1 U4797 ( .A(N1388), .B(n7202), .Y(n7050) );
  INVX1 U4798 ( .A(n5161), .Y(n7202) );
  NAND3X1 U4799 ( .A(n7205), .B(n5461), .C(N2880), .Y(n5161) );
  INVX1 U4800 ( .A(N2777), .Y(n5461) );
  INVX1 U4801 ( .A(n6480), .Y(n7205) );
  NAND2X1 U4802 ( .A(n4612), .B(n4298), .Y(n6480) );
  INVX1 U4803 ( .A(N3336), .Y(n4298) );
  NOR2X1 U4804 ( .A(n4297), .B(n4080), .Y(n4612) );
  INVX1 U4805 ( .A(n4128), .Y(n4080) );
  OAI21X1 U4806 ( .A(n3477), .B(n4070), .C(n7051), .Y(n4128) );
  AOI22X1 U4807 ( .A(n7052), .B(n7053), .C(Gy[31]), .D(n7054), .Y(n7051) );
  OAI21X1 U4808 ( .A(n3546), .B(n3547), .C(n3481), .Y(n7054) );
  NAND2X1 U4809 ( .A(n4293), .B(n4131), .Y(n3552) );
  NAND2X1 U4810 ( .A(IntSignal[1]), .B(n3540), .Y(n3547) );
  INVX1 U4811 ( .A(IntSignal[0]), .Y(n3540) );
  NOR2X1 U4812 ( .A(\regX[6][5] ), .B(n7055), .Y(n7053) );
  NAND2X1 U4813 ( .A(n3848), .B(n3849), .Y(n7055) );
  INVX1 U4814 ( .A(\regX[6][7] ), .Y(n3849) );
  INVX1 U4815 ( .A(\regX[6][6] ), .Y(n3848) );
  NOR2X1 U4816 ( .A(n4297), .B(n7056), .Y(n7052) );
  OAI21X1 U4817 ( .A(n7057), .B(n7058), .C(n3846), .Y(n7056) );
  INVX1 U4818 ( .A(\regX[6][4] ), .Y(n3846) );
  NAND2X1 U4819 ( .A(\regX[6][3] ), .B(\regX[6][2] ), .Y(n7058) );
  NAND2X1 U4820 ( .A(\regX[6][1] ), .B(\regX[6][0] ), .Y(n7057) );
  INVX1 U4821 ( .A(fGx[31]), .Y(n4070) );
  INVX1 U4822 ( .A(n3546), .Y(n4131) );
  NAND3X1 U4823 ( .A(n7059), .B(n7060), .C(OPMode[0]), .Y(n3546) );
  INVX1 U4824 ( .A(OPMode[1]), .Y(n7059) );
  INVX1 U4825 ( .A(n5725), .Y(n5457) );
  NAND2X1 U4826 ( .A(IntSignal[1]), .B(IntSignal[0]), .Y(n5725) );
  NAND3X1 U4827 ( .A(n4293), .B(OPMode[0]), .C(n4256), .Y(n4297) );
  INVX1 U4828 ( .A(dx[0]), .Y(n7004) );
  NAND3X1 U4829 ( .A(n7246), .B(n3864), .C(N2777), .Y(n3943) );
  INVX1 U4830 ( .A(N2549), .Y(n3864) );
  NAND3X1 U4831 ( .A(n4293), .B(n4250), .C(n4256), .Y(n5827) );
  INVX1 U4832 ( .A(n3549), .Y(n4256) );
  NAND2X1 U4833 ( .A(OPMode[1]), .B(n7060), .Y(n3549) );
  INVX1 U4834 ( .A(OPMode[2]), .Y(n7060) );
  INVX1 U4835 ( .A(OPMode[0]), .Y(n4250) );
  INVX1 U4836 ( .A(n5453), .Y(n4293) );
  NAND2X1 U4837 ( .A(IntSignal[0]), .B(n3554), .Y(n5453) );
  INVX1 U4838 ( .A(IntSignal[1]), .Y(n3554) );
  AND2X1 U4839 ( .A(N3194), .B(bCE), .Y(\U3/U100/Z_6 ) );
  NOR2X1 U4840 ( .A(n7061), .B(n7062), .Y(N1582) );
  OR2X1 U4841 ( .A(n7063), .B(n7064), .Y(n7062) );
  INVX1 U4842 ( .A(N1776), .Y(n7061) );
  XOR2X1 U4843 ( .A(N1776), .B(n7065), .Y(N1581) );
  NOR2X1 U4844 ( .A(n7064), .B(n7063), .Y(n7065) );
  XOR2X1 U4845 ( .A(n7063), .B(n7064), .Y(N1580) );
  NAND3X1 U4846 ( .A(N1773), .B(n7066), .C(N1774), .Y(n7064) );
  INVX1 U4847 ( .A(N1775), .Y(n7063) );
  XOR2X1 U4848 ( .A(N1774), .B(n7067), .Y(N1579) );
  AND2X1 U4849 ( .A(n7066), .B(N1773), .Y(n7067) );
  XOR2X1 U4850 ( .A(N1773), .B(n7066), .Y(N1578) );
  OAI21X1 U4851 ( .A(n7068), .B(n3764), .C(n7069), .Y(n7066) );
  OAI21X1 U4852 ( .A(N1742), .B(n7070), .C(N1772), .Y(n7069) );
  XOR2X1 U4853 ( .A(n7071), .B(n7068), .Y(N1577) );
  INVX1 U4854 ( .A(n7070), .Y(n7068) );
  OAI21X1 U4855 ( .A(n7072), .B(n3763), .C(n7073), .Y(n7070) );
  OAI21X1 U4856 ( .A(N1741), .B(n7074), .C(N1771), .Y(n7073) );
  XOR2X1 U4857 ( .A(N1772), .B(n3764), .Y(n7071) );
  INVX1 U4858 ( .A(N1742), .Y(n3764) );
  XOR2X1 U4859 ( .A(n7075), .B(n7072), .Y(N1576) );
  INVX1 U4860 ( .A(n7074), .Y(n7072) );
  OAI21X1 U4861 ( .A(n7076), .B(n3762), .C(n7077), .Y(n7074) );
  OAI21X1 U4862 ( .A(N1740), .B(n7078), .C(N1770), .Y(n7077) );
  XOR2X1 U4863 ( .A(N1771), .B(n3763), .Y(n7075) );
  INVX1 U4864 ( .A(N1741), .Y(n3763) );
  XOR2X1 U4865 ( .A(n7079), .B(n7076), .Y(N1575) );
  INVX1 U4866 ( .A(n7078), .Y(n7076) );
  OAI21X1 U4867 ( .A(n7080), .B(n3761), .C(n7081), .Y(n7078) );
  OAI21X1 U4868 ( .A(N1739), .B(n7082), .C(N1769), .Y(n7081) );
  XOR2X1 U4869 ( .A(N1770), .B(n3762), .Y(n7079) );
  INVX1 U4870 ( .A(N1740), .Y(n3762) );
  XOR2X1 U4871 ( .A(n7083), .B(n7080), .Y(N1574) );
  INVX1 U4872 ( .A(n7082), .Y(n7080) );
  OAI21X1 U4873 ( .A(n7084), .B(n3760), .C(n7085), .Y(n7082) );
  OAI21X1 U4874 ( .A(N1738), .B(n7086), .C(N1768), .Y(n7085) );
  XOR2X1 U4875 ( .A(N1769), .B(n3761), .Y(n7083) );
  INVX1 U4876 ( .A(N1739), .Y(n3761) );
  XOR2X1 U4877 ( .A(n7087), .B(n7084), .Y(N1573) );
  INVX1 U4878 ( .A(n7086), .Y(n7084) );
  OAI21X1 U4879 ( .A(n3759), .B(n7088), .C(n7089), .Y(n7086) );
  OAI21X1 U4880 ( .A(n7090), .B(N1737), .C(N1767), .Y(n7089) );
  INVX1 U4881 ( .A(n7088), .Y(n7090) );
  XOR2X1 U4882 ( .A(N1768), .B(n3760), .Y(n7087) );
  INVX1 U4883 ( .A(N1738), .Y(n3760) );
  XOR2X1 U4884 ( .A(n7088), .B(n7091), .Y(N1572) );
  XOR2X1 U4885 ( .A(N1767), .B(n3759), .Y(n7091) );
  INVX1 U4886 ( .A(N1737), .Y(n3759) );
  OAI21X1 U4887 ( .A(N1736), .B(n7092), .C(n7093), .Y(n7088) );
  OAI21X1 U4888 ( .A(n3758), .B(n7094), .C(n7095), .Y(n7093) );
  INVX1 U4889 ( .A(N1736), .Y(n3758) );
  INVX1 U4890 ( .A(n7094), .Y(n7092) );
  XOR2X1 U4891 ( .A(n7094), .B(n7096), .Y(N1571) );
  XOR2X1 U4892 ( .A(n7095), .B(N1736), .Y(n7096) );
  INVX1 U4893 ( .A(N1766), .Y(n7095) );
  NAND2X1 U4894 ( .A(N1765), .B(N1735), .Y(n7094) );
  XOR2X1 U4895 ( .A(N1765), .B(N1735), .Y(N1570) );
  NOR2X1 U4896 ( .A(n7097), .B(n7098), .Y(N1552) );
  NAND2X1 U4897 ( .A(N1715), .B(n7099), .Y(n7098) );
  INVX1 U4898 ( .A(N1716), .Y(n7097) );
  XOR2X1 U4899 ( .A(N1716), .B(n7100), .Y(N1551) );
  AND2X1 U4900 ( .A(n7099), .B(N1715), .Y(n7100) );
  XOR2X1 U4901 ( .A(N1715), .B(n7099), .Y(N1550) );
  OAI21X1 U4902 ( .A(n7101), .B(n3784), .C(n7102), .Y(n7099) );
  OAI21X1 U4903 ( .A(N1684), .B(n7103), .C(N1714), .Y(n7102) );
  XOR2X1 U4904 ( .A(n7104), .B(n7101), .Y(N1549) );
  INVX1 U4905 ( .A(n7103), .Y(n7101) );
  OAI21X1 U4906 ( .A(n7105), .B(n3783), .C(n7106), .Y(n7103) );
  OAI21X1 U4907 ( .A(N1683), .B(n7107), .C(N1713), .Y(n7106) );
  XOR2X1 U4908 ( .A(N1714), .B(n3784), .Y(n7104) );
  INVX1 U4909 ( .A(N1684), .Y(n3784) );
  XOR2X1 U4910 ( .A(n7108), .B(n7105), .Y(N1548) );
  INVX1 U4911 ( .A(n7107), .Y(n7105) );
  OAI21X1 U4912 ( .A(n7109), .B(n3782), .C(n7110), .Y(n7107) );
  OAI21X1 U4913 ( .A(N1682), .B(n7111), .C(N1712), .Y(n7110) );
  XOR2X1 U4914 ( .A(N1713), .B(n3783), .Y(n7108) );
  INVX1 U4915 ( .A(N1683), .Y(n3783) );
  XOR2X1 U4916 ( .A(n7112), .B(n7109), .Y(N1547) );
  INVX1 U4917 ( .A(n7111), .Y(n7109) );
  OAI21X1 U4918 ( .A(n7113), .B(n3781), .C(n7114), .Y(n7111) );
  OAI21X1 U4919 ( .A(N1681), .B(n7115), .C(N1711), .Y(n7114) );
  XOR2X1 U4920 ( .A(N1712), .B(n3782), .Y(n7112) );
  INVX1 U4921 ( .A(N1682), .Y(n3782) );
  XOR2X1 U4922 ( .A(n7116), .B(n7113), .Y(N1546) );
  INVX1 U4923 ( .A(n7115), .Y(n7113) );
  OAI21X1 U4924 ( .A(n7117), .B(n3780), .C(n7118), .Y(n7115) );
  OAI21X1 U4925 ( .A(N1680), .B(n7119), .C(N1710), .Y(n7118) );
  XOR2X1 U4926 ( .A(N1711), .B(n3781), .Y(n7116) );
  INVX1 U4927 ( .A(N1681), .Y(n3781) );
  XOR2X1 U4928 ( .A(n7120), .B(n7117), .Y(N1545) );
  INVX1 U4929 ( .A(n7119), .Y(n7117) );
  OAI21X1 U4930 ( .A(n3779), .B(n7121), .C(n7122), .Y(n7119) );
  OAI21X1 U4931 ( .A(n7123), .B(N1679), .C(N1709), .Y(n7122) );
  INVX1 U4932 ( .A(n7121), .Y(n7123) );
  XOR2X1 U4933 ( .A(N1710), .B(n3780), .Y(n7120) );
  INVX1 U4934 ( .A(N1680), .Y(n3780) );
  XOR2X1 U4935 ( .A(n7121), .B(n7124), .Y(N1544) );
  XOR2X1 U4936 ( .A(N1709), .B(n3779), .Y(n7124) );
  INVX1 U4937 ( .A(N1679), .Y(n3779) );
  OAI21X1 U4938 ( .A(N1678), .B(n7125), .C(n7126), .Y(n7121) );
  OAI21X1 U4939 ( .A(n3778), .B(n7127), .C(n7128), .Y(n7126) );
  INVX1 U4940 ( .A(N1678), .Y(n3778) );
  INVX1 U4941 ( .A(n7127), .Y(n7125) );
  XOR2X1 U4942 ( .A(n7127), .B(n7129), .Y(N1543) );
  XOR2X1 U4943 ( .A(n7128), .B(N1678), .Y(n7129) );
  INVX1 U4944 ( .A(N1708), .Y(n7128) );
  NAND2X1 U4945 ( .A(N1707), .B(N1677), .Y(n7127) );
  XOR2X1 U4946 ( .A(N1707), .B(N1677), .Y(N1542) );
  NOR2X1 U4947 ( .A(n7130), .B(n7131), .Y(N1522) );
  OR2X1 U4948 ( .A(n7132), .B(n7133), .Y(n7131) );
  INVX1 U4949 ( .A(N1656), .Y(n7130) );
  XOR2X1 U4950 ( .A(N1656), .B(n7134), .Y(N1521) );
  NOR2X1 U4951 ( .A(n7133), .B(n7132), .Y(n7134) );
  XOR2X1 U4952 ( .A(n7132), .B(n7133), .Y(N1520) );
  NAND3X1 U4953 ( .A(N1653), .B(n7135), .C(N1654), .Y(n7133) );
  INVX1 U4954 ( .A(N1655), .Y(n7132) );
  XOR2X1 U4955 ( .A(N1654), .B(n7136), .Y(N1519) );
  AND2X1 U4956 ( .A(n7135), .B(N1653), .Y(n7136) );
  XOR2X1 U4957 ( .A(N1653), .B(n7135), .Y(N1518) );
  OAI21X1 U4958 ( .A(n7137), .B(n3803), .C(n7138), .Y(n7135) );
  OAI21X1 U4959 ( .A(N1622), .B(n7139), .C(N1652), .Y(n7138) );
  XOR2X1 U4960 ( .A(n7140), .B(n7137), .Y(N1517) );
  INVX1 U4961 ( .A(n7139), .Y(n7137) );
  OAI21X1 U4962 ( .A(n7141), .B(n3802), .C(n7142), .Y(n7139) );
  OAI21X1 U4963 ( .A(N1621), .B(n7143), .C(N1651), .Y(n7142) );
  XOR2X1 U4964 ( .A(N1652), .B(n3803), .Y(n7140) );
  INVX1 U4965 ( .A(N1622), .Y(n3803) );
  XOR2X1 U4966 ( .A(n7144), .B(n7141), .Y(N1516) );
  INVX1 U4967 ( .A(n7143), .Y(n7141) );
  OAI21X1 U4968 ( .A(n7145), .B(n3801), .C(n7146), .Y(n7143) );
  OAI21X1 U4969 ( .A(N1620), .B(n7147), .C(N1650), .Y(n7146) );
  XOR2X1 U4970 ( .A(N1651), .B(n3802), .Y(n7144) );
  INVX1 U4971 ( .A(N1621), .Y(n3802) );
  XOR2X1 U4972 ( .A(n7148), .B(n7145), .Y(N1515) );
  INVX1 U4973 ( .A(n7147), .Y(n7145) );
  OAI21X1 U4974 ( .A(n7149), .B(n3800), .C(n7150), .Y(n7147) );
  OAI21X1 U4975 ( .A(N1619), .B(n7151), .C(N1649), .Y(n7150) );
  XOR2X1 U4976 ( .A(N1650), .B(n3801), .Y(n7148) );
  INVX1 U4977 ( .A(N1620), .Y(n3801) );
  XOR2X1 U4978 ( .A(n7152), .B(n7149), .Y(N1514) );
  INVX1 U4979 ( .A(n7151), .Y(n7149) );
  OAI21X1 U4980 ( .A(n7153), .B(n3799), .C(n7154), .Y(n7151) );
  OAI21X1 U4981 ( .A(N1618), .B(n7155), .C(N1648), .Y(n7154) );
  XOR2X1 U4982 ( .A(N1649), .B(n3800), .Y(n7152) );
  INVX1 U4983 ( .A(N1619), .Y(n3800) );
  XOR2X1 U4984 ( .A(n7156), .B(n7153), .Y(N1513) );
  INVX1 U4985 ( .A(n7155), .Y(n7153) );
  OAI21X1 U4986 ( .A(n3798), .B(n7157), .C(n7158), .Y(n7155) );
  OAI21X1 U4987 ( .A(n7159), .B(N1617), .C(N1647), .Y(n7158) );
  INVX1 U4988 ( .A(n7157), .Y(n7159) );
  XOR2X1 U4989 ( .A(N1648), .B(n3799), .Y(n7156) );
  INVX1 U4990 ( .A(N1618), .Y(n3799) );
  XOR2X1 U4991 ( .A(n7157), .B(n7160), .Y(N1512) );
  XOR2X1 U4992 ( .A(N1647), .B(n3798), .Y(n7160) );
  INVX1 U4993 ( .A(N1617), .Y(n3798) );
  OAI21X1 U4994 ( .A(N1616), .B(n7161), .C(n7162), .Y(n7157) );
  OAI21X1 U4995 ( .A(n3797), .B(n7163), .C(n7164), .Y(n7162) );
  INVX1 U4996 ( .A(N1616), .Y(n3797) );
  INVX1 U4997 ( .A(n7163), .Y(n7161) );
  XOR2X1 U4998 ( .A(n7163), .B(n7165), .Y(N1511) );
  XOR2X1 U4999 ( .A(n7164), .B(N1616), .Y(n7165) );
  INVX1 U5000 ( .A(N1646), .Y(n7164) );
  NAND2X1 U5001 ( .A(N1645), .B(N1615), .Y(n7163) );
  XOR2X1 U5002 ( .A(N1645), .B(N1615), .Y(N1510) );
  XOR2X1 U5003 ( .A(N1417), .B(n7166), .Y(N1402) );
  AND2X1 U5004 ( .A(n7167), .B(N1416), .Y(n7166) );
  XOR2X1 U5005 ( .A(N1416), .B(n7167), .Y(N1401) );
  NOR2X1 U5006 ( .A(n7168), .B(n7169), .Y(n7167) );
  XOR2X1 U5007 ( .A(n7168), .B(n7169), .Y(N1400) );
  NAND3X1 U5008 ( .A(N1413), .B(n7170), .C(N1414), .Y(n7169) );
  INVX1 U5009 ( .A(N1415), .Y(n7168) );
  XNOR2X1 U5010 ( .A(N1414), .B(n7171), .Y(N1399) );
  NAND2X1 U5011 ( .A(N1413), .B(n7170), .Y(n7171) );
  XOR2X1 U5012 ( .A(n7170), .B(N1413), .Y(N1398) );
  OAI21X1 U5013 ( .A(n7172), .B(n3911), .C(n7173), .Y(n7170) );
  OAI21X1 U5014 ( .A(N1382), .B(n7174), .C(N1412), .Y(n7173) );
  INVX1 U5015 ( .A(N1382), .Y(n3911) );
  INVX1 U5016 ( .A(n7174), .Y(n7172) );
  XOR2X1 U5017 ( .A(n7174), .B(n7175), .Y(N1397) );
  XOR2X1 U5018 ( .A(N1412), .B(N1382), .Y(n7175) );
  OAI21X1 U5019 ( .A(n7176), .B(n3910), .C(n7177), .Y(n7174) );
  OAI21X1 U5020 ( .A(N1381), .B(n7178), .C(N1411), .Y(n7177) );
  XOR2X1 U5021 ( .A(n7179), .B(n7176), .Y(N1396) );
  INVX1 U5022 ( .A(n7178), .Y(n7176) );
  OAI21X1 U5023 ( .A(n7180), .B(n3909), .C(n7181), .Y(n7178) );
  OAI21X1 U5024 ( .A(N1380), .B(n7182), .C(N1410), .Y(n7181) );
  XOR2X1 U5025 ( .A(N1411), .B(n3910), .Y(n7179) );
  INVX1 U5026 ( .A(N1381), .Y(n3910) );
  XOR2X1 U5027 ( .A(n7183), .B(n7180), .Y(N1395) );
  INVX1 U5028 ( .A(n7182), .Y(n7180) );
  OAI21X1 U5029 ( .A(n7184), .B(n3908), .C(n7185), .Y(n7182) );
  OAI21X1 U5030 ( .A(N1379), .B(n7186), .C(N1409), .Y(n7185) );
  XOR2X1 U5031 ( .A(N1410), .B(n3909), .Y(n7183) );
  INVX1 U5032 ( .A(N1380), .Y(n3909) );
  XOR2X1 U5033 ( .A(n7187), .B(n7184), .Y(N1394) );
  INVX1 U5034 ( .A(n7186), .Y(n7184) );
  OAI21X1 U5035 ( .A(n7188), .B(n3907), .C(n7189), .Y(n7186) );
  OAI21X1 U5036 ( .A(N1378), .B(n7190), .C(N1408), .Y(n7189) );
  XOR2X1 U5037 ( .A(N1409), .B(n3908), .Y(n7187) );
  INVX1 U5038 ( .A(N1379), .Y(n3908) );
  XOR2X1 U5039 ( .A(n7191), .B(n7188), .Y(N1393) );
  INVX1 U5040 ( .A(n7190), .Y(n7188) );
  OAI21X1 U5041 ( .A(n7192), .B(n3906), .C(n7193), .Y(n7190) );
  OAI21X1 U5042 ( .A(N1377), .B(n7194), .C(N3443), .Y(n7193) );
  INVX1 U5043 ( .A(N1377), .Y(n3906) );
  XOR2X1 U5044 ( .A(N1408), .B(n3907), .Y(n7191) );
  INVX1 U5045 ( .A(N1378), .Y(n3907) );
  XOR2X1 U5046 ( .A(n7195), .B(n7192), .Y(N1392) );
  INVX1 U5047 ( .A(n7194), .Y(n7192) );
  OAI21X1 U5048 ( .A(n7048), .B(n3905), .C(n7196), .Y(n7194) );
  NAND3X1 U5049 ( .A(N3441), .B(n7197), .C(N1375), .Y(n7196) );
  XOR2X1 U5050 ( .A(n7040), .B(N1377), .Y(n7195) );
  INVX1 U5051 ( .A(N3443), .Y(n7040) );
  XOR2X1 U5052 ( .A(n7198), .B(n7199), .Y(N1391) );
  NAND2X1 U5053 ( .A(N1375), .B(N3441), .Y(n7199) );
  OAI21X1 U5054 ( .A(n7048), .B(n3905), .C(n7197), .Y(n7198) );
  NAND2X1 U5055 ( .A(n7048), .B(n3905), .Y(n7197) );
  INVX1 U5056 ( .A(N1376), .Y(n3905) );
  INVX1 U5057 ( .A(N3442), .Y(n7048) );
  XOR2X1 U5058 ( .A(N3441), .B(N1375), .Y(N1390) );
endmodule


module WRAP_CANNY ( DataBus, AddressBus, ControlBus, AddrRegRow, AddrRegCol, 
        bWE, bCE, InDataToCanny, OutDataFromCanny, OPMode, bOPEnable, dReadReg, 
        dWriteReg, Breq, Bgnt, clk, bReset );
  inout [7:0] DataBus;
  inout [31:0] AddressBus;
  output [2:0] AddrRegRow;
  output [2:0] AddrRegCol;
  output [7:0] InDataToCanny;
  input [7:0] OutDataFromCanny;
  output [2:0] OPMode;
  output [3:0] dReadReg;
  output [3:0] dWriteReg;
  input Bgnt, clk, bReset;
  output bWE, bCE, bOPEnable, Breq;
  inout ControlBus;
  wire   IntEnable, n47, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n54, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134;
  tri   [7:0] DataBus;
  tri   [31:0] AddressBus;
  tri   AddressBus_7;
  tri   AddressBus_6;
  tri   AddressBus_5;
  tri   AddressBus_4;
  tri   AddressBus_3;
  tri   AddressBus_2;
  tri   AddressBus_1;
  tri   AddressBus_0;
  tri   ControlBus;
  tri   [7:0] OutDataFromCanny;
  tran( AddressBus_7, AddressBus[7]);
  tran( AddressBus_6, AddressBus[6]);
  tran( AddressBus_5, AddressBus[5]);
  tran( AddressBus_4, AddressBus[4]);
  tran( AddressBus_3, AddressBus[3]);
  tran( AddressBus_2, AddressBus[2]);
  tran( AddressBus_1, AddressBus[1]);
  tran( AddressBus_0, AddressBus[0]);

  DFFPOSX1 IntEnable_reg ( .D(n84), .CLK(clk), .Q(IntEnable) );
  DFFPOSX1 \InDataToCanny_reg[0]  ( .D(n83), .CLK(clk), .Q(InDataToCanny[0])
         );
  DFFPOSX1 \InDataToCanny_reg[2]  ( .D(n81), .CLK(clk), .Q(InDataToCanny[2])
         );
  DFFPOSX1 \InDataToCanny_reg[4]  ( .D(n79), .CLK(clk), .Q(InDataToCanny[4])
         );
  DFFPOSX1 \InDataToCanny_reg[6]  ( .D(n77), .CLK(clk), .Q(InDataToCanny[6])
         );
  DFFPOSX1 \InDataToCanny_reg[7]  ( .D(n76), .CLK(clk), .Q(InDataToCanny[7])
         );
  DFFPOSX1 \InDataToCanny_reg[5]  ( .D(n78), .CLK(clk), .Q(InDataToCanny[5])
         );
  DFFPOSX1 \InDataToCanny_reg[3]  ( .D(n80), .CLK(clk), .Q(InDataToCanny[3])
         );
  DFFPOSX1 \InDataToCanny_reg[1]  ( .D(n82), .CLK(clk), .Q(InDataToCanny[1])
         );
  DFFPOSX1 \dWriteReg_reg[3]  ( .D(n56), .CLK(clk), .Q(dWriteReg[3]) );
  DFFPOSX1 \dWriteReg_reg[2]  ( .D(n57), .CLK(clk), .Q(dWriteReg[2]) );
  DFFPOSX1 \dWriteReg_reg[1]  ( .D(n58), .CLK(clk), .Q(dWriteReg[1]) );
  DFFPOSX1 \dWriteReg_reg[0]  ( .D(n59), .CLK(clk), .Q(dWriteReg[0]) );
  DFFPOSX1 \dReadReg_reg[3]  ( .D(n60), .CLK(clk), .Q(dReadReg[3]) );
  DFFPOSX1 \dReadReg_reg[2]  ( .D(n61), .CLK(clk), .Q(dReadReg[2]) );
  DFFPOSX1 \dReadReg_reg[1]  ( .D(n62), .CLK(clk), .Q(dReadReg[1]) );
  DFFPOSX1 \dReadReg_reg[0]  ( .D(n63), .CLK(clk), .Q(dReadReg[0]) );
  DFFPOSX1 bOPEnable_reg ( .D(n64), .CLK(clk), .Q(bOPEnable) );
  DFFPOSX1 \OPMode_reg[2]  ( .D(n65), .CLK(clk), .Q(OPMode[2]) );
  DFFPOSX1 \OPMode_reg[1]  ( .D(n66), .CLK(clk), .Q(OPMode[1]) );
  DFFPOSX1 \OPMode_reg[0]  ( .D(n67), .CLK(clk), .Q(OPMode[0]) );
  DFFPOSX1 bCE_reg ( .D(n68), .CLK(clk), .Q(bCE) );
  DFFPOSX1 bWE_reg ( .D(n69), .CLK(clk), .Q(bWE) );
  DFFPOSX1 \AddrRegCol_reg[2]  ( .D(n70), .CLK(clk), .Q(AddrRegCol[2]) );
  DFFPOSX1 \AddrRegCol_reg[1]  ( .D(n71), .CLK(clk), .Q(AddrRegCol[1]) );
  DFFPOSX1 \AddrRegCol_reg[0]  ( .D(n72), .CLK(clk), .Q(AddrRegCol[0]) );
  DFFPOSX1 \AddrRegRow_reg[2]  ( .D(n73), .CLK(clk), .Q(AddrRegRow[2]) );
  DFFPOSX1 \AddrRegRow_reg[1]  ( .D(n74), .CLK(clk), .Q(AddrRegRow[1]) );
  DFFPOSX1 \AddrRegRow_reg[0]  ( .D(n75), .CLK(clk), .Q(AddrRegRow[0]) );
  DFFPOSX1 Breq_reg ( .D(n55), .CLK(clk), .Q(Breq) );
  TBUFX1 \DataBus_tri[0]  ( .A(n134), .EN(n47), .Y(DataBus[0]) );
  TBUFX1 \DataBus_tri[1]  ( .A(n133), .EN(n47), .Y(DataBus[1]) );
  TBUFX1 \DataBus_tri[2]  ( .A(n132), .EN(n47), .Y(DataBus[2]) );
  TBUFX1 \DataBus_tri[3]  ( .A(n131), .EN(n47), .Y(DataBus[3]) );
  TBUFX1 \DataBus_tri[4]  ( .A(n130), .EN(n47), .Y(DataBus[4]) );
  TBUFX1 \DataBus_tri[5]  ( .A(n129), .EN(n47), .Y(DataBus[5]) );
  TBUFX1 \DataBus_tri[6]  ( .A(n128), .EN(n47), .Y(DataBus[6]) );
  TBUFX1 \DataBus_tri[7]  ( .A(n127), .EN(n47), .Y(DataBus[7]) );
  TBUFX1 ControlBus_tri ( .A(1'b1), .EN(IntEnable), .Y(ControlBus) );
  INVX1 U3 ( .A(OutDataFromCanny[7]), .Y(n127) );
  INVX1 U4 ( .A(OutDataFromCanny[6]), .Y(n128) );
  INVX1 U5 ( .A(OutDataFromCanny[5]), .Y(n129) );
  INVX1 U6 ( .A(OutDataFromCanny[4]), .Y(n130) );
  INVX1 U7 ( .A(OutDataFromCanny[3]), .Y(n131) );
  INVX1 U8 ( .A(OutDataFromCanny[2]), .Y(n132) );
  INVX1 U9 ( .A(OutDataFromCanny[1]), .Y(n133) );
  INVX1 U10 ( .A(OutDataFromCanny[0]), .Y(n134) );
  AND2X1 U11 ( .A(bReset), .B(n54), .Y(n84) );
  OAI21X1 U12 ( .A(IntEnable), .B(n85), .C(n86), .Y(n54) );
  INVX1 U13 ( .A(Bgnt), .Y(n85) );
  INVX1 U14 ( .A(n87), .Y(n83) );
  MUX2X1 U15 ( .B(DataBus[0]), .A(InDataToCanny[0]), .S(n88), .Y(n87) );
  INVX1 U16 ( .A(n89), .Y(n82) );
  MUX2X1 U17 ( .B(DataBus[1]), .A(InDataToCanny[1]), .S(n88), .Y(n89) );
  INVX1 U18 ( .A(n90), .Y(n81) );
  MUX2X1 U19 ( .B(DataBus[2]), .A(InDataToCanny[2]), .S(n88), .Y(n90) );
  INVX1 U20 ( .A(n91), .Y(n80) );
  MUX2X1 U21 ( .B(DataBus[3]), .A(InDataToCanny[3]), .S(n88), .Y(n91) );
  INVX1 U22 ( .A(n92), .Y(n79) );
  MUX2X1 U23 ( .B(DataBus[4]), .A(InDataToCanny[4]), .S(n88), .Y(n92) );
  INVX1 U24 ( .A(n93), .Y(n78) );
  MUX2X1 U25 ( .B(DataBus[5]), .A(InDataToCanny[5]), .S(n88), .Y(n93) );
  INVX1 U26 ( .A(n94), .Y(n77) );
  MUX2X1 U27 ( .B(DataBus[6]), .A(InDataToCanny[6]), .S(n88), .Y(n94) );
  INVX1 U28 ( .A(n95), .Y(n76) );
  MUX2X1 U29 ( .B(DataBus[7]), .A(InDataToCanny[7]), .S(n88), .Y(n95) );
  NAND3X1 U30 ( .A(n96), .B(n97), .C(n98), .Y(n88) );
  INVX1 U31 ( .A(n99), .Y(n75) );
  MUX2X1 U32 ( .B(AddressBus_5), .A(AddrRegRow[0]), .S(n86), .Y(n99) );
  INVX1 U33 ( .A(n100), .Y(n74) );
  MUX2X1 U34 ( .B(AddressBus_6), .A(AddrRegRow[1]), .S(n86), .Y(n100) );
  INVX1 U35 ( .A(n101), .Y(n73) );
  MUX2X1 U36 ( .B(AddressBus_7), .A(AddrRegRow[2]), .S(n86), .Y(n101) );
  INVX1 U37 ( .A(n102), .Y(n72) );
  MUX2X1 U38 ( .B(AddressBus_2), .A(AddrRegCol[0]), .S(n86), .Y(n102) );
  INVX1 U39 ( .A(n103), .Y(n71) );
  MUX2X1 U40 ( .B(AddressBus_3), .A(AddrRegCol[1]), .S(n86), .Y(n103) );
  INVX1 U41 ( .A(n104), .Y(n70) );
  MUX2X1 U42 ( .B(AddressBus_4), .A(AddrRegCol[2]), .S(n86), .Y(n104) );
  INVX1 U43 ( .A(n105), .Y(n69) );
  MUX2X1 U44 ( .B(AddressBus_1), .A(bWE), .S(n86), .Y(n105) );
  INVX1 U45 ( .A(n106), .Y(n68) );
  MUX2X1 U46 ( .B(AddressBus_0), .A(bCE), .S(n86), .Y(n106) );
  INVX1 U47 ( .A(n107), .Y(n67) );
  MUX2X1 U48 ( .B(AddressBus[24]), .A(OPMode[0]), .S(n86), .Y(n107) );
  INVX1 U49 ( .A(n108), .Y(n66) );
  MUX2X1 U50 ( .B(AddressBus[25]), .A(OPMode[1]), .S(n86), .Y(n108) );
  INVX1 U51 ( .A(n109), .Y(n65) );
  MUX2X1 U52 ( .B(AddressBus[26]), .A(OPMode[2]), .S(n86), .Y(n109) );
  INVX1 U53 ( .A(n110), .Y(n64) );
  MUX2X1 U54 ( .B(AddressBus[27]), .A(bOPEnable), .S(n86), .Y(n110) );
  INVX1 U55 ( .A(n111), .Y(n63) );
  MUX2X1 U56 ( .B(AddressBus[16]), .A(dReadReg[0]), .S(n86), .Y(n111) );
  INVX1 U57 ( .A(n112), .Y(n62) );
  MUX2X1 U58 ( .B(AddressBus[17]), .A(dReadReg[1]), .S(n86), .Y(n112) );
  INVX1 U59 ( .A(n113), .Y(n61) );
  MUX2X1 U60 ( .B(AddressBus[18]), .A(dReadReg[2]), .S(n86), .Y(n113) );
  INVX1 U61 ( .A(n114), .Y(n60) );
  MUX2X1 U62 ( .B(AddressBus[19]), .A(dReadReg[3]), .S(n86), .Y(n114) );
  INVX1 U63 ( .A(n115), .Y(n59) );
  MUX2X1 U64 ( .B(AddressBus[20]), .A(dWriteReg[0]), .S(n86), .Y(n115) );
  INVX1 U65 ( .A(n116), .Y(n58) );
  MUX2X1 U66 ( .B(AddressBus[21]), .A(dWriteReg[1]), .S(n86), .Y(n116) );
  INVX1 U67 ( .A(n117), .Y(n57) );
  MUX2X1 U68 ( .B(AddressBus[22]), .A(dWriteReg[2]), .S(n86), .Y(n117) );
  INVX1 U69 ( .A(n118), .Y(n56) );
  MUX2X1 U70 ( .B(AddressBus[23]), .A(dWriteReg[3]), .S(n86), .Y(n118) );
  NOR2X1 U71 ( .A(n119), .B(n120), .Y(n55) );
  INVX1 U72 ( .A(bReset), .Y(n120) );
  AOI22X1 U73 ( .A(n121), .B(n122), .C(Breq), .D(n98), .Y(n119) );
  NOR2X1 U74 ( .A(IntEnable), .B(Bgnt), .Y(n121) );
  NOR2X1 U75 ( .A(n97), .B(n123), .Y(n47) );
  NAND2X1 U76 ( .A(n98), .B(n96), .Y(n123) );
  INVX1 U77 ( .A(AddressBus_0), .Y(n96) );
  INVX1 U78 ( .A(n86), .Y(n98) );
  NAND2X1 U79 ( .A(IntEnable), .B(n122), .Y(n86) );
  INVX1 U80 ( .A(n124), .Y(n122) );
  NAND3X1 U81 ( .A(AddressBus[30]), .B(n125), .C(n126), .Y(n124) );
  NOR2X1 U82 ( .A(AddressBus[31]), .B(AddressBus[29]), .Y(n126) );
  INVX1 U83 ( .A(AddressBus[28]), .Y(n125) );
  INVX1 U84 ( .A(AddressBus_1), .Y(n97) );
endmodule


module Arbiter ( BREQn, BGNTn );
  input [3:0] BREQn;
  output [3:0] BGNTn;
  wire   BREQn_3, \BREQn[2] , n7, n8, n9, n10, n11, n12;
  assign BREQn_3 = BREQn[3];
  assign BGNTn[2] = \BREQn[2] ;
  assign \BREQn[2]  = BREQn[2];

  NOR2X1 U1 ( .A(n7), .B(n8), .Y(BGNTn[3]) );
  NAND2X1 U2 ( .A(BREQn_3), .B(n9), .Y(n8) );
  NAND2X1 U3 ( .A(n10), .B(n11), .Y(n7) );
  NOR2X1 U4 ( .A(n10), .B(n12), .Y(BGNTn[1]) );
  NAND2X1 U5 ( .A(n9), .B(n11), .Y(n12) );
  INVX1 U6 ( .A(\BREQn[2] ), .Y(n11) );
  INVX1 U7 ( .A(BREQn[1]), .Y(n10) );
  NOR2X1 U8 ( .A(\BREQn[2] ), .B(n9), .Y(BGNTn[0]) );
  INVX1 U9 ( .A(BREQn[0]), .Y(n9) );
endmodule


module systemtop ( Serial_out, clk, Breq, Bgnt, DataBus, AddressBus, 
        ControlBus, bReset );
  inout [7:0] DataBus;
  inout [31:0] AddressBus;
  input clk, Breq, bReset;
  output Serial_out, Bgnt;
  inout ControlBus;
  wire   Breqn_3, Bgntn_3, bCE, bWE, Load_XMT_datareg, Byte_ready, T_byte,
         Canny_bWE, Canny_bCE, bOPEnable;
  wire   [1:0] Breqn;
  wire   [1:0] Bgntn;
  wire   [7:0] InData;
  wire   [7:0] OutData;
  wire   [17:0] Address;
  wire   [7:0] DataToUART;
  wire   [2:0] AddrRegRow;
  wire   [2:0] AddrRegCol;
  wire   [7:0] DataToCanny;
  wire   [2:0] OPMode;
  wire   [3:0] dReadReg;
  wire   [3:0] dWriteReg;
  tri   Serial_out;
  tri   [7:0] DataBus;
  tri   [31:0] AddressBus;
  tri   ControlBus;
  tri   [7:0] DataFromCanny;

  SRAM SRAM_01 ( .InData(InData), .OutData(OutData), .Address(Address), .bCE(
        bCE), .bWE(bWE) );
  WRAP_SRAM WRAP_SRAM_01 ( .DataBus(DataBus), .AddressBus(AddressBus), 
        .ControlBus(ControlBus), .InData(InData), .OutData(OutData), .Address(
        Address), .bCE(bCE), .bWE(bWE), .Breq(Breqn[0]), .Bgnt(Bgntn[0]), 
        .clk(clk), .bReset(bReset) );
  UART_XMTR UART_XMTR_01 ( .Serial_out(Serial_out), .Data_Bus(DataToUART), 
        .Load_XMT_datareg(Load_XMT_datareg), .Byte_ready(Byte_ready), .T_byte(
        T_byte), .Clock(clk), .rst_b(bReset) );
  WRAP_UART WRAP_UART_01 ( .DataBus(DataBus), .AddressBus(AddressBus), 
        .ControlBus(ControlBus), .InData(DataToUART), .Load_XMT_datareg(
        Load_XMT_datareg), .Byte_ready(Byte_ready), .T_byte(T_byte), .Breq(
        Breqn[1]), .Bgnt(Bgntn[1]), .clk(clk), .bReset(bReset) );
  CannyEdge CannyEdge_01 ( .dAddrRegRow(AddrRegRow), .dAddrRegCol(AddrRegCol), 
        .bWE(Canny_bWE), .bCE(Canny_bCE), .InData(DataToCanny), .OutData(
        DataFromCanny), .OPMode(OPMode), .bOPEnable(bOPEnable), .dReadReg(
        dReadReg), .dWriteReg(dWriteReg), .clk(clk), .rst_b(bReset) );
  WRAP_CANNY WRAP_CANNY_01 ( .DataBus(DataBus), .AddressBus(AddressBus), 
        .ControlBus(ControlBus), .AddrRegRow(AddrRegRow), .AddrRegCol(
        AddrRegCol), .bWE(Canny_bWE), .bCE(Canny_bCE), .InDataToCanny(
        DataToCanny), .OutDataFromCanny(DataFromCanny), .OPMode(OPMode), 
        .bOPEnable(bOPEnable), .dReadReg(dReadReg), .dWriteReg(dWriteReg), 
        .Breq(Breqn_3), .Bgnt(Bgntn_3), .clk(clk), .bReset(bReset) );
  Arbiter Arbiter_01 ( .BREQn({Breqn_3, Breq, Breqn}), .BGNTn({Bgntn_3, Bgnt, 
        Bgntn}) );
endmodule

